module Instruction_decode(clk, ireset, irq, inst, c, z, read_strobe,
     write_strobe, interrupt_ack, next_interrupt_enabled,
     interrupt_enabled, zsel, csel, wsel, pcsel, stsel, werf, wesp);
  input clk, ireset, irq, c, z, interrupt_enabled;
  input [17:0] inst;
  output read_strobe, write_strobe, interrupt_ack,
       next_interrupt_enabled, werf, wesp;
  output [2:0] zsel, csel, wsel;
  output [1:0] pcsel, stsel;

  wire AA_111, AA_117, AA_125, AA_129, AA_136, AA_139, AA_147, AA_148, AA_150, AA_153, 
       AA_154, AA_162, AA_164, AA_165, AA_167, AA_168, AA_169, AA_170, AA_171, AA_173, 
       AA_176, AA_178, AA_179, AA_180, AA_181, AA_182, AA_191, AA_207, AA_214, AA_215, 
       AA_217, AA_220, AA_223, AA_224, AA_225, AA_226, AA_227, AA_228, AA_229, AA_230, 
       AA_231, AA_232, AA_241, AA_242, AA_245, AA_253, AA_260, AA_262, AA_263, AA_264, 
       AA_269, AA_27, AA_272, AA_273, AA_274, AA_275, AA_279, AA_280, AA_281, AA_282, 
       AA_283, AA_284, AA_285, AA_292, AA_294, AA_298, AA_302, AA_308, AA_311, AA_313, 
       AA_325, AA_326, AA_328, AA_334, AA_335, AA_336, AA_340, AA_341, AA_342, AA_372, 
       AA_386, AA_391, AA_392, AA_393, AA_394, AA_395, AA_396, AA_397, AA_398, AA_399, 
       AA_400, AA_401, AA_402, AA_403, AA_404, AA_405, AA_406, AA_407, AA_408, AA_409, 
       AA_410, AA_411, AA_416, AA_419, AA_420, AA_421, AA_422, AA_423, AA_424, AA_425, 
       AA_426, AA_427, AA_428, AA_429, AA_430, AA_431, AA_432, AA_433, AA_434, AA_435, 
       AA_436, AA_441, AA_442, AA_443, AA_444, AA_445, AA_446, AA_447, AA_448, AA_449, 
       AA_450, AA_451, AA_452, AA_453, AA_454, AA_455, AA_456, AA_458, AA_459, AA_460, 
       AA_461, AA_462, AA_463, AA_464, AA_53, AA_79, AA_83, AA_93, BB_0_30, BB_0_3021, 
       BB_0_30211, BB_0_31, BB_0_311, BB_0_3110, BB_0_31100, BB_0_3121, BB_0_320, BB_0_321, BB_0_3211, BB_100_30, 
       BB_100_30222221, BB_100_31, BB_100_310, BB_100_3101, BB_100_31011, BB_100_310221, BB_100_311, BB_100_3110, BB_100_31101, BB_100_311011, 
       BB_100_3111, BB_100_31110, BB_100_31111, BB_100_311111, BB_100_31120, BB_100_31121, BB_100_311211, BB_100_3121, BB_100_31211, BB_100_312110, 
       BB_100_3222220, BB_100_32222201, BB_100_3222221, BB_100_32222211, BB_13_30, BB_13_300, BB_13_3000, BB_13_301, BB_13_3011, BB_13_3021, 
       BB_13_31, BB_13_310, BB_13_320, BB_183_31, BB_183_310, BB_183_3101, BB_183_31011, BB_183_310221, BB_183_311, BB_183_3110, 
       BB_183_31101, BB_183_311011, BB_183_3110111, BB_183_3111, BB_183_31110, BB_183_31111, BB_183_311111, BB_183_3111111, BB_183_31111110, BB_183_311111100, 
       BB_183_31120, BB_183_311201, BB_183_31121, BB_183_311211, BB_183_3112111, BB_183_3121, BB_183_31211, BB_183_312111, BB_183_3121111, BB_233_31, 
       BB_233_310, BB_233_3101, BB_233_31011, BB_233_310221, BB_233_311, BB_233_3110, BB_233_31101, BB_233_311011, BB_233_3111, BB_233_31110, 
       BB_233_31111, BB_233_311111, BB_233_31120, BB_233_31121, BB_233_311211, BB_233_3121, BB_233_31211, BB_286_30, BB_286_30222221, BB_286_31, 
       BB_286_310, BB_286_3101, BB_286_31011, BB_286_310221, BB_286_311, BB_286_3110, BB_286_31101, BB_286_311011, BB_286_3111, BB_286_31110, 
       BB_286_31111, BB_286_311111, BB_286_31120, BB_286_31121, BB_286_311211, BB_286_3121, BB_286_31211, BB_286_312110, BB_286_3222220, BB_286_32222201, 
       BB_286_3222221, BB_286_32222211, BB_28_30, BB_28_301, BB_28_3010, BB_28_31, BB_28_311, BB_28_3111, BB_28_321, BB_28_3211, 
       BB_28_32111, BB_343_31, BB_343_310, BB_343_3100, BB_343_311, BB_343_3121, BB_343_31211, BB_350_30, BB_350_301, BB_350_3010, 
       BB_350_31, BB_350_311, BB_350_321, BB_360_31, BB_361_30, BB_361_301, BB_361_3011, BB_361_30110, BB_361_301100, BB_361_31, 
       BB_361_310, BB_361_3101, BB_361_31010, BB_361_31011, BB_361_311, BB_361_3111, BB_361_31110, BB_361_3120, BB_361_3121, BB_361_31211, 
       BB_361_312110, BB_361_312120, BB_361_3121201, BB_361_321, BB_361_3211, BB_361_32110, BB_361_321100, BB_361_32111, BB_373_30, BB_373_300, 
       BB_373_3000, BB_373_30000, BB_373_31, BB_373_310, BB_373_31020, BB_373_311, BB_373_321, BB_387_31, BB_40_30, BB_40_300, 
       BB_40_31, BB_40_310, BB_40_311, BB_40_3111, BB_40_3121, BB_40_320, BB_40_3201, BB_40_32010, BB_40_32021, BB_40_321, 
       BB_40_3211, BB_40_321220, BB_40_3221, BB_61_30, BB_61_300, BB_61_3000, BB_61_30000, BB_61_31, BB_61_310, BB_61_3101, 
       BB_61_311, BB_61_3110, BB_61_3120, BB_61_320, BB_61_3201, BB_61_32010, BB_61_321, BB_61_3210, BB_61_3211, BB_61_32110, 
       BB_61_321100, BB_61_3220, BB_61_3221, BB_84_30, BB_84_300, BB_84_3000, BB_84_301, BB_84_3010, BB_84_3011, BB_84_31, 
       BB_84_310, BB_84_3101, BB_84_311, BB_84_3111, BB_84_31121, BB_84_320, BB_84_321, BB_84_3210, BB_84_3211, BB_97_30, 
       BB_97_31, BB_97_311, BB_99_31, csel[0], csel[1], csel[2], interrupt_ack, next_interrupt_enabled, pcsel[0], pcsel[1], 
       read_strobe, stsel[0], stsel[1], werf, wesp, write_strobe, wsel[0], wsel[1], zsel[0], zsel[1], zsel[2];

NEMR4T g1(.s(zsel[0]), .d(BB_0_30), .b(vdd), .g(inst[14]));
NEMR4T g2(.s(BB_0_30), .d(AA_463), .b(vdd), .g(inst[16]));
NEMR4T g3(.s(AA_463), .d(AA_458), .b(vdd), .g(inst[13]));
NEMR4T g4(.s(AA_458), .d(AA_441), .b(vdd), .g(irq));
NEMR4T g5(.s(AA_441), .d(AA_391), .b(gnd), .g(inst[17]));
NEMR4T g6(.s(AA_391), .d(vdd), .b(vdd), .g(inst[15]));
NEMR4T g7(.s(AA_458), .d(AA_442), .b(vdd), .g(inst[17]));
NEMR4T g8(.s(AA_442), .d(AA_392), .b(vdd), .g(ireset));
NEMR4T g9(.s(AA_392), .d(gnd), .b(gnd), .g(vdd));
NEMR4T g10(.s(AA_442), .d(AA_393), .b(gnd), .g(ireset));
NEMR4T g11(.s(AA_393), .d(vdd), .b(gnd), .g(vdd));
NEMR4T g12(.s(BB_0_30), .d(AA_443), .b(gnd), .g(inst[16]));
NEMR4T g13(.s(AA_443), .d(AA_396), .b(vdd), .g(irq));
NEMR4T g14(.s(AA_396), .d(AA_394), .b(vdd), .g(inst[17]));
NEMR4T g15(.s(AA_394), .d(vdd), .b(gnd), .g(inst[15]));
NEMR4T g16(.s(AA_396), .d(AA_395), .b(vdd), .g(ireset));
NEMR4T g17(.s(AA_395), .d(gnd), .b(vdd), .g(inst[15]));
NEMR4T g18(.s(AA_396), .d(AA_391), .b(gnd), .g(ireset));
NEMR4T g19(.s(BB_0_30), .d(AA_444), .b(vdd), .g(inst[13]));
NEMR4T g20(.s(AA_444), .d(AA_398), .b(gnd), .g(inst[17]));
NEMR4T g21(.s(AA_398), .d(AA_397), .b(vdd), .g(ireset));
NEMR4T g22(.s(AA_397), .d(gnd), .b(gnd), .g(inst[15]));
NEMR4T g23(.s(AA_398), .d(AA_394), .b(gnd), .g(ireset));
NEMR4T g24(.s(BB_0_30), .d(BB_0_3021), .b(gnd), .g(inst[13]));
NEMR4T g25(.s(BB_0_3021), .d(BB_0_30211), .b(gnd), .g(irq));
NEMR4T g26(.s(BB_0_30211), .d(AA_442), .b(vdd), .g(inst[17]));
NEMR4T g27(.s(BB_0_30211), .d(AA_398), .b(gnd), .g(inst[17]));
NEMR4T g28(.s(BB_0_30), .d(AA_445), .b(gnd), .g(irq));
NEMR4T g29(.s(AA_445), .d(AA_399), .b(gnd), .g(inst[17]));
NEMR4T g30(.s(AA_399), .d(AA_395), .b(vdd), .g(ireset));
NEMR4T g31(.s(AA_399), .d(AA_391), .b(gnd), .g(ireset));
NEMR4T g32(.s(zsel[0]), .d(BB_0_31), .b(gnd), .g(inst[14]));
NEMR4T g33(.s(BB_0_31), .d(AA_446), .b(vdd), .g(inst[16]));
NEMR4T g34(.s(AA_446), .d(AA_442), .b(vdd), .g(inst[13]));
NEMR4T g35(.s(BB_0_31), .d(BB_0_311), .b(gnd), .g(inst[16]));
NEMR4T g36(.s(BB_0_311), .d(BB_0_3110), .b(vdd), .g(inst[13]));
NEMR4T g37(.s(BB_0_3110), .d(BB_0_31100), .b(vdd), .g(irq));
NEMR4T g38(.s(BB_0_31100), .d(AA_393), .b(vdd), .g(inst[17]));
NEMR4T g39(.s(BB_0_3110), .d(AA_442), .b(gnd), .g(inst[17]));
NEMR4T g40(.s(BB_0_311), .d(AA_443), .b(gnd), .g(inst[13]));
NEMR4T g41(.s(BB_0_31), .d(BB_0_3121), .b(gnd), .g(inst[13]));
NEMR4T g42(.s(BB_0_3121), .d(AA_442), .b(gnd), .g(irq));
NEMR4T g43(.s(zsel[0]), .d(BB_0_320), .b(vdd), .g(inst[16]));
NEMR4T g44(.s(BB_0_320), .d(AA_447), .b(gnd), .g(inst[13]));
NEMR4T g45(.s(AA_447), .d(AA_442), .b(vdd), .g(irq));
NEMR4T g46(.s(zsel[0]), .d(BB_0_321), .b(gnd), .g(inst[16]));
NEMR4T g47(.s(BB_0_321), .d(AA_459), .b(vdd), .g(inst[13]));
NEMR4T g48(.s(AA_459), .d(AA_448), .b(gnd), .g(irq));
NEMR4T g49(.s(AA_448), .d(AA_442), .b(vdd), .g(inst[17]));
NEMR4T g50(.s(BB_0_321), .d(BB_0_3211), .b(gnd), .g(inst[13]));
NEMR4T g51(.s(BB_0_3211), .d(AA_444), .b(vdd), .g(irq));
NEMR4T g52(.s(zsel[1]), .d(BB_13_30), .b(vdd), .g(inst[14]));
NEMR4T g53(.s(BB_13_30), .d(BB_13_300), .b(vdd), .g(inst[16]));
NEMR4T g54(.s(BB_13_300), .d(BB_13_3000), .b(vdd), .g(inst[13]));
NEMR4T g55(.s(BB_13_3000), .d(AA_449), .b(vdd), .g(irq));
NEMR4T g56(.s(AA_449), .d(AA_400), .b(gnd), .g(inst[17]));
NEMR4T g57(.s(AA_400), .d(AA_391), .b(vdd), .g(ireset));
NEMR4T g58(.s(AA_400), .d(gnd), .b(gnd), .g(inst[15]));
NEMR4T g59(.s(BB_13_3000), .d(AA_392), .b(vdd), .g(inst[17]));
NEMR4T g60(.s(BB_13_300), .d(AA_450), .b(gnd), .g(irq));
NEMR4T g61(.s(AA_450), .d(AA_401), .b(gnd), .g(inst[17]));
NEMR4T g62(.s(AA_401), .d(AA_392), .b(vdd), .g(ireset));
NEMR4T g63(.s(BB_13_30), .d(BB_13_301), .b(gnd), .g(inst[16]));
NEMR4T g64(.s(BB_13_301), .d(BB_13_3011), .b(gnd), .g(inst[13]));
NEMR4T g65(.s(BB_13_3011), .d(AA_402), .b(vdd), .g(irq));
NEMR4T g66(.s(AA_402), .d(AA_400), .b(vdd), .g(inst[17]));
NEMR4T g67(.s(AA_402), .d(AA_395), .b(gnd), .g(ireset));
NEMR4T g68(.s(BB_13_3011), .d(AA_403), .b(gnd), .g(inst[17]));
NEMR4T g69(.s(AA_403), .d(AA_397), .b(gnd), .g(ireset));
NEMR4T g70(.s(BB_13_30), .d(BB_13_3021), .b(gnd), .g(inst[13]));
NEMR4T g71(.s(BB_13_3021), .d(AA_450), .b(vdd), .g(irq));
NEMR4T g72(.s(BB_13_3021), .d(AA_404), .b(gnd), .g(irq));
NEMR4T g73(.s(AA_404), .d(AA_392), .b(vdd), .g(inst[17]));
NEMR4T g74(.s(zsel[1]), .d(BB_13_31), .b(gnd), .g(inst[14]));
NEMR4T g75(.s(BB_13_31), .d(BB_13_310), .b(vdd), .g(inst[16]));
NEMR4T g76(.s(BB_13_310), .d(AA_27), .b(vdd), .g(inst[13]));
NEMR4T g77(.s(AA_27), .d(AA_406), .b(vdd), .g(irq));
NEMR4T g78(.s(AA_406), .d(AA_405), .b(vdd), .g(inst[17]));
NEMR4T g79(.s(AA_405), .d(AA_394), .b(vdd), .g(ireset));
NEMR4T g80(.s(AA_405), .d(gnd), .b(vdd), .g(inst[15]));
NEMR4T g81(.s(AA_406), .d(AA_397), .b(gnd), .g(ireset));
NEMR4T g82(.s(BB_13_310), .d(AA_404), .b(gnd), .g(irq));
NEMR4T g83(.s(BB_13_310), .d(AA_401), .b(gnd), .g(inst[17]));
NEMR4T g84(.s(BB_13_31), .d(AA_460), .b(gnd), .g(inst[16]));
NEMR4T g85(.s(AA_460), .d(AA_451), .b(gnd), .g(inst[13]));
NEMR4T g86(.s(AA_451), .d(AA_392), .b(vdd), .g(irq));
NEMR4T g87(.s(AA_451), .d(AA_407), .b(gnd), .g(irq));
NEMR4T g88(.s(AA_407), .d(AA_392), .b(vdd), .g(inst[17]));
NEMR4T g89(.s(AA_407), .d(AA_403), .b(gnd), .g(inst[17]));
NEMR4T g90(.s(zsel[1]), .d(BB_13_320), .b(vdd), .g(inst[16]));
NEMR4T g91(.s(BB_13_320), .d(AA_27), .b(gnd), .g(inst[13]));
NEMR4T g92(.s(BB_13_320), .d(AA_408), .b(gnd), .g(irq));
NEMR4T g93(.s(AA_408), .d(AA_403), .b(gnd), .g(inst[17]));
NEMR4T g94(.s(BB_13_320), .d(AA_409), .b(gnd), .g(inst[17]));
NEMR4T g95(.s(AA_409), .d(AA_395), .b(gnd), .g(ireset));
NEMR4T g96(.s(zsel[1]), .d(AA_464), .b(gnd), .g(inst[16]));
NEMR4T g97(.s(AA_464), .d(AA_392), .b(vdd), .g(inst[13]));
NEMR4T g98(.s(AA_464), .d(AA_461), .b(gnd), .g(inst[13]));
NEMR4T g99(.s(AA_461), .d(AA_452), .b(gnd), .g(irq));
NEMR4T g100(.s(AA_452), .d(AA_410), .b(gnd), .g(inst[17]));
NEMR4T g101(.s(AA_410), .d(AA_392), .b(vdd), .g(ireset));
NEMR4T g102(.s(AA_410), .d(AA_395), .b(gnd), .g(ireset));
NEMR4T g103(.s(zsel[2]), .d(BB_28_30), .b(vdd), .g(inst[14]));
NEMR4T g104(.s(BB_28_30), .d(BB_28_301), .b(gnd), .g(inst[16]));
NEMR4T g105(.s(BB_28_301), .d(BB_28_3010), .b(vdd), .g(inst[13]));
NEMR4T g106(.s(BB_28_3010), .d(AA_411), .b(vdd), .g(irq));
NEMR4T g107(.s(AA_411), .d(AA_394), .b(gnd), .g(inst[17]));
NEMR4T g108(.s(BB_28_3010), .d(AA_442), .b(vdd), .g(inst[17]));
NEMR4T g109(.s(BB_28_3010), .d(AA_399), .b(gnd), .g(inst[17]));
NEMR4T g110(.s(BB_28_301), .d(AA_444), .b(gnd), .g(irq));
NEMR4T g111(.s(zsel[2]), .d(BB_28_31), .b(gnd), .g(inst[14]));
NEMR4T g112(.s(BB_28_31), .d(BB_28_311), .b(gnd), .g(inst[16]));
NEMR4T g113(.s(BB_28_311), .d(AA_442), .b(vdd), .g(inst[13]));
NEMR4T g114(.s(BB_28_311), .d(BB_28_3111), .b(gnd), .g(inst[13]));
NEMR4T g115(.s(BB_28_3111), .d(AA_444), .b(gnd), .g(irq));
NEMR4T g116(.s(zsel[2]), .d(AA_442), .b(vdd), .g(inst[16]));
NEMR4T g117(.s(zsel[2]), .d(BB_28_321), .b(gnd), .g(inst[16]));
NEMR4T g118(.s(BB_28_321), .d(BB_28_3211), .b(gnd), .g(inst[13]));
NEMR4T g119(.s(BB_28_3211), .d(AA_442), .b(vdd), .g(irq));
NEMR4T g120(.s(BB_28_3211), .d(BB_28_32111), .b(gnd), .g(irq));
NEMR4T g121(.s(BB_28_32111), .d(AA_442), .b(vdd), .g(inst[17]));
NEMR4T g122(.s(BB_28_32111), .d(AA_399), .b(gnd), .g(inst[17]));
NEMR4T g123(.s(csel[0]), .d(BB_40_30), .b(vdd), .g(inst[3]));
NEMR4T g124(.s(BB_40_30), .d(BB_40_300), .b(vdd), .g(inst[14]));
NEMR4T g125(.s(BB_40_300), .d(AA_446), .b(vdd), .g(inst[16]));
NEMR4T g126(.s(BB_40_300), .d(AA_416), .b(gnd), .g(inst[13]));
NEMR4T g127(.s(AA_416), .d(AA_445), .b(gnd), .g(irq));
NEMR4T g128(.s(AA_416), .d(AA_398), .b(gnd), .g(inst[17]));
NEMR4T g129(.s(BB_40_30), .d(AA_416), .b(gnd), .g(inst[14]));
NEMR4T g130(.s(csel[0]), .d(BB_40_31), .b(gnd), .g(inst[3]));
NEMR4T g131(.s(BB_40_31), .d(BB_40_310), .b(vdd), .g(inst[14]));
NEMR4T g132(.s(BB_40_310), .d(AA_463), .b(vdd), .g(inst[16]));
NEMR4T g133(.s(BB_40_31), .d(BB_40_311), .b(gnd), .g(inst[14]));
NEMR4T g134(.s(BB_40_311), .d(BB_40_3111), .b(gnd), .g(inst[16]));
NEMR4T g135(.s(BB_40_3111), .d(AA_416), .b(vdd), .g(inst[13]));
NEMR4T g136(.s(BB_40_31), .d(AA_416), .b(vdd), .g(inst[16]));
NEMR4T g137(.s(BB_40_31), .d(BB_40_3121), .b(gnd), .g(inst[16]));
NEMR4T g138(.s(BB_40_3121), .d(AA_416), .b(gnd), .g(inst[13]));
NEMR4T g139(.s(csel[0]), .d(BB_40_320), .b(vdd), .g(inst[14]));
NEMR4T g140(.s(BB_40_320), .d(BB_40_3201), .b(gnd), .g(inst[16]));
NEMR4T g141(.s(BB_40_3201), .d(BB_40_32010), .b(vdd), .g(inst[13]));
NEMR4T g142(.s(BB_40_32010), .d(AA_394), .b(vdd), .g(irq));
NEMR4T g143(.s(BB_40_32010), .d(AA_442), .b(gnd), .g(irq));
NEMR4T g144(.s(BB_40_320), .d(BB_40_32021), .b(gnd), .g(inst[13]));
NEMR4T g145(.s(BB_40_32021), .d(AA_396), .b(vdd), .g(irq));
NEMR4T g146(.s(BB_40_32021), .d(AA_448), .b(gnd), .g(irq));
NEMR4T g147(.s(csel[0]), .d(BB_40_321), .b(gnd), .g(inst[14]));
NEMR4T g148(.s(BB_40_321), .d(AA_53), .b(vdd), .g(inst[16]));
NEMR4T g149(.s(AA_53), .d(AA_399), .b(vdd), .g(irq));
NEMR4T g150(.s(BB_40_321), .d(BB_40_3211), .b(gnd), .g(inst[16]));
NEMR4T g151(.s(BB_40_3211), .d(AA_53), .b(gnd), .g(inst[13]));
NEMR4T g152(.s(BB_40_321), .d(BB_40_321220), .b(vdd), .g(irq));
NEMR4T g153(.s(BB_40_321220), .d(AA_394), .b(vdd), .g(inst[17]));
NEMR4T g154(.s(BB_40_321), .d(AA_448), .b(gnd), .g(irq));
NEMR4T g155(.s(csel[0]), .d(BB_40_3221), .b(gnd), .g(inst[16]));
NEMR4T g156(.s(BB_40_3221), .d(AA_53), .b(vdd), .g(inst[13]));
NEMR4T g157(.s(csel[1]), .d(BB_61_30), .b(vdd), .g(inst[3]));
NEMR4T g158(.s(BB_61_30), .d(BB_61_300), .b(vdd), .g(inst[14]));
NEMR4T g159(.s(BB_61_300), .d(BB_61_3000), .b(vdd), .g(inst[16]));
NEMR4T g160(.s(BB_61_3000), .d(BB_61_30000), .b(vdd), .g(inst[13]));
NEMR4T g161(.s(BB_61_30000), .d(AA_441), .b(vdd), .g(irq));
NEMR4T g162(.s(BB_61_300), .d(AA_448), .b(vdd), .g(inst[13]));
NEMR4T g163(.s(BB_61_30), .d(AA_416), .b(vdd), .g(inst[16]));
NEMR4T g164(.s(BB_61_30), .d(AA_83), .b(gnd), .g(inst[16]));
NEMR4T g165(.s(AA_83), .d(AA_79), .b(gnd), .g(inst[13]));
NEMR4T g166(.s(AA_79), .d(AA_445), .b(gnd), .g(irq));
NEMR4T g167(.s(csel[1]), .d(BB_61_31), .b(gnd), .g(inst[3]));
NEMR4T g168(.s(BB_61_31), .d(BB_61_310), .b(vdd), .g(inst[14]));
NEMR4T g169(.s(BB_61_310), .d(AA_446), .b(vdd), .g(inst[16]));
NEMR4T g170(.s(BB_61_310), .d(BB_61_3101), .b(gnd), .g(inst[16]));
NEMR4T g171(.s(BB_61_3101), .d(AA_448), .b(vdd), .g(inst[13]));
NEMR4T g172(.s(BB_61_310), .d(AA_79), .b(gnd), .g(inst[13]));
NEMR4T g173(.s(BB_61_31), .d(BB_61_311), .b(gnd), .g(inst[14]));
NEMR4T g174(.s(BB_61_311), .d(BB_61_3110), .b(vdd), .g(inst[16]));
NEMR4T g175(.s(BB_61_3110), .d(AA_444), .b(vdd), .g(inst[13]));
NEMR4T g176(.s(BB_61_3110), .d(AA_445), .b(gnd), .g(irq));
NEMR4T g177(.s(BB_61_311), .d(AA_83), .b(gnd), .g(inst[16]));
NEMR4T g178(.s(BB_61_31), .d(BB_61_3120), .b(vdd), .g(inst[16]));
NEMR4T g179(.s(BB_61_3120), .d(AA_444), .b(gnd), .g(inst[13]));
NEMR4T g180(.s(csel[1]), .d(BB_61_320), .b(vdd), .g(inst[14]));
NEMR4T g181(.s(BB_61_320), .d(BB_61_3201), .b(gnd), .g(inst[16]));
NEMR4T g182(.s(BB_61_3201), .d(BB_61_32010), .b(vdd), .g(inst[13]));
NEMR4T g183(.s(BB_61_32010), .d(AA_411), .b(vdd), .g(irq));
NEMR4T g184(.s(BB_61_320), .d(AA_459), .b(gnd), .g(inst[13]));
NEMR4T g185(.s(csel[1]), .d(BB_61_321), .b(gnd), .g(inst[14]));
NEMR4T g186(.s(BB_61_321), .d(BB_61_3210), .b(vdd), .g(inst[16]));
NEMR4T g187(.s(BB_61_3210), .d(AA_443), .b(vdd), .g(inst[13]));
NEMR4T g188(.s(BB_61_321), .d(BB_61_3211), .b(gnd), .g(inst[16]));
NEMR4T g189(.s(BB_61_3211), .d(BB_61_32110), .b(vdd), .g(inst[13]));
NEMR4T g190(.s(BB_61_32110), .d(BB_61_321100), .b(vdd), .g(irq));
NEMR4T g191(.s(BB_61_321100), .d(AA_391), .b(vdd), .g(inst[17]));
NEMR4T g192(.s(BB_61_321100), .d(AA_397), .b(vdd), .g(ireset));
NEMR4T g193(.s(BB_61_321100), .d(AA_394), .b(gnd), .g(ireset));
NEMR4T g194(.s(BB_61_321), .d(AA_448), .b(gnd), .g(irq));
NEMR4T g195(.s(csel[1]), .d(BB_61_3220), .b(vdd), .g(inst[16]));
NEMR4T g196(.s(BB_61_3220), .d(AA_443), .b(gnd), .g(inst[13]));
NEMR4T g197(.s(csel[1]), .d(BB_61_3221), .b(gnd), .g(inst[16]));
NEMR4T g198(.s(BB_61_3221), .d(AA_445), .b(vdd), .g(inst[13]));
NEMR4T g199(.s(BB_61_3221), .d(AA_447), .b(gnd), .g(inst[13]));
NEMR4T g200(.s(BB_61_3221), .d(AA_444), .b(gnd), .g(irq));
NEMR4T g201(.s(csel[2]), .d(BB_84_30), .b(vdd), .g(inst[14]));
NEMR4T g202(.s(BB_84_30), .d(BB_84_300), .b(vdd), .g(inst[16]));
NEMR4T g203(.s(BB_84_300), .d(BB_84_3000), .b(vdd), .g(inst[13]));
NEMR4T g204(.s(BB_84_3000), .d(AA_449), .b(vdd), .g(irq));
NEMR4T g205(.s(BB_84_3000), .d(AA_409), .b(gnd), .g(inst[17]));
NEMR4T g206(.s(BB_84_300), .d(AA_408), .b(gnd), .g(irq));
NEMR4T g207(.s(BB_84_30), .d(BB_84_301), .b(gnd), .g(inst[16]));
NEMR4T g208(.s(BB_84_301), .d(BB_84_3010), .b(vdd), .g(inst[13]));
NEMR4T g209(.s(BB_84_3010), .d(AA_419), .b(vdd), .g(irq));
NEMR4T g210(.s(AA_419), .d(AA_405), .b(gnd), .g(inst[17]));
NEMR4T g211(.s(BB_84_301), .d(BB_84_3011), .b(gnd), .g(inst[13]));
NEMR4T g212(.s(BB_84_3011), .d(AA_402), .b(vdd), .g(irq));
NEMR4T g213(.s(BB_84_301), .d(AA_403), .b(gnd), .g(inst[17]));
NEMR4T g214(.s(BB_84_30), .d(AA_404), .b(vdd), .g(inst[13]));
NEMR4T g215(.s(BB_84_30), .d(AA_453), .b(gnd), .g(inst[13]));
NEMR4T g216(.s(AA_453), .d(AA_420), .b(gnd), .g(irq));
NEMR4T g217(.s(AA_420), .d(AA_392), .b(vdd), .g(inst[17]));
NEMR4T g218(.s(AA_420), .d(AA_409), .b(gnd), .g(inst[17]));
NEMR4T g219(.s(BB_84_30), .d(AA_450), .b(gnd), .g(irq));
NEMR4T g220(.s(csel[2]), .d(BB_84_31), .b(gnd), .g(inst[14]));
NEMR4T g221(.s(BB_84_31), .d(BB_84_310), .b(vdd), .g(inst[16]));
NEMR4T g222(.s(BB_84_310), .d(AA_392), .b(vdd), .g(inst[13]));
NEMR4T g223(.s(BB_84_310), .d(BB_84_3101), .b(gnd), .g(inst[13]));
NEMR4T g224(.s(BB_84_3101), .d(AA_392), .b(gnd), .g(irq));
NEMR4T g225(.s(BB_84_31), .d(BB_84_311), .b(gnd), .g(inst[16]));
NEMR4T g226(.s(BB_84_311), .d(AA_421), .b(vdd), .g(inst[13]));
NEMR4T g227(.s(AA_421), .d(AA_392), .b(vdd), .g(irq));
NEMR4T g228(.s(BB_84_311), .d(BB_84_3111), .b(gnd), .g(inst[13]));
NEMR4T g229(.s(BB_84_3111), .d(AA_454), .b(vdd), .g(irq));
NEMR4T g230(.s(AA_454), .d(AA_392), .b(vdd), .g(inst[17]));
NEMR4T g231(.s(AA_454), .d(AA_422), .b(gnd), .g(inst[17]));
NEMR4T g232(.s(AA_422), .d(AA_392), .b(gnd), .g(ireset));
NEMR4T g233(.s(BB_84_3111), .d(AA_93), .b(gnd), .g(irq));
NEMR4T g234(.s(AA_93), .d(AA_409), .b(gnd), .g(inst[17]));
NEMR4T g235(.s(BB_84_311), .d(BB_84_31121), .b(gnd), .g(irq));
NEMR4T g236(.s(BB_84_31121), .d(AA_392), .b(vdd), .g(inst[17]));
NEMR4T g237(.s(BB_84_31121), .d(AA_423), .b(gnd), .g(inst[17]));
NEMR4T g238(.s(AA_423), .d(AA_392), .b(vdd), .g(ireset));
NEMR4T g239(.s(AA_423), .d(AA_397), .b(gnd), .g(ireset));
NEMR4T g240(.s(csel[2]), .d(BB_84_320), .b(vdd), .g(inst[16]));
NEMR4T g241(.s(BB_84_320), .d(AA_421), .b(gnd), .g(inst[13]));
NEMR4T g242(.s(csel[2]), .d(BB_84_321), .b(gnd), .g(inst[16]));
NEMR4T g243(.s(BB_84_321), .d(BB_84_3210), .b(vdd), .g(inst[13]));
NEMR4T g244(.s(BB_84_3210), .d(AA_93), .b(gnd), .g(irq));
NEMR4T g245(.s(BB_84_321), .d(BB_84_3211), .b(gnd), .g(inst[13]));
NEMR4T g246(.s(BB_84_3211), .d(AA_450), .b(vdd), .g(irq));
NEMR4T g247(.s(wsel[0]), .d(BB_97_30), .b(vdd), .g(inst[14]));
NEMR4T g248(.s(BB_97_30), .d(AA_392), .b(vdd), .g(inst[17]));
NEMR4T g249(.s(BB_97_30), .d(AA_393), .b(gnd), .g(inst[17]));
NEMR4T g250(.s(wsel[0]), .d(BB_97_31), .b(gnd), .g(inst[14]));
NEMR4T g251(.s(BB_97_31), .d(AA_391), .b(vdd), .g(inst[13]));
NEMR4T g252(.s(BB_97_31), .d(BB_97_311), .b(gnd), .g(inst[13]));
NEMR4T g253(.s(BB_97_311), .d(AA_395), .b(vdd), .g(inst[17]));
NEMR4T g254(.s(BB_97_311), .d(AA_391), .b(gnd), .g(inst[17]));
NEMR4T g255(.s(BB_97_31), .d(AA_397), .b(vdd), .g(inst[17]));
NEMR4T g256(.s(BB_97_31), .d(AA_394), .b(gnd), .g(inst[17]));
NEMR4T g257(.s(wsel[1]), .d(AA_392), .b(vdd), .g(inst[14]));
NEMR4T g258(.s(wsel[1]), .d(BB_99_31), .b(gnd), .g(inst[14]));
NEMR4T g259(.s(BB_99_31), .d(vdd), .b(vdd), .g(inst[15]));
NEMR4T g260(.s(BB_99_31), .d(gnd), .b(gnd), .g(inst[15]));
NEMR4T g261(.s(pcsel[1]), .d(BB_100_30), .b(vdd), .g(inst[12]));
NEMR4T g262(.s(BB_100_30), .d(AA_179), .b(vdd), .g(inst[14]));
NEMR4T g263(.s(AA_179), .d(AA_178), .b(vdd), .g(inst[16]));
NEMR4T g264(.s(AA_178), .d(AA_167), .b(gnd), .g(inst[13]));
NEMR4T g265(.s(AA_167), .d(AA_411), .b(vdd), .g(irq));
NEMR4T g266(.s(AA_167), .d(AA_424), .b(gnd), .g(irq));
NEMR4T g267(.s(AA_424), .d(AA_393), .b(vdd), .g(ireset));
NEMR4T g268(.s(AA_167), .d(AA_425), .b(vdd), .g(inst[17]));
NEMR4T g269(.s(AA_425), .d(AA_393), .b(gnd), .g(ireset));
NEMR4T g270(.s(AA_167), .d(AA_426), .b(gnd), .g(inst[17]));
NEMR4T g271(.s(AA_426), .d(AA_391), .b(gnd), .g(ireset));
NEMR4T g272(.s(AA_179), .d(AA_169), .b(gnd), .g(inst[13]));
NEMR4T g273(.s(AA_169), .d(AA_168), .b(vdd), .g(irq));
NEMR4T g274(.s(AA_168), .d(AA_401), .b(vdd), .g(inst[17]));
NEMR4T g275(.s(AA_168), .d(AA_427), .b(gnd), .g(inst[17]));
NEMR4T g276(.s(AA_427), .d(AA_395), .b(vdd), .g(ireset));
NEMR4T g277(.s(AA_169), .d(AA_147), .b(gnd), .g(irq));
NEMR4T g278(.s(AA_147), .d(AA_428), .b(gnd), .g(inst[17]));
NEMR4T g279(.s(AA_428), .d(AA_394), .b(gnd), .g(ireset));
NEMR4T g280(.s(BB_100_30), .d(AA_182), .b(gnd), .g(inst[14]));
NEMR4T g281(.s(AA_182), .d(AA_148), .b(vdd), .g(inst[16]));
NEMR4T g282(.s(AA_148), .d(AA_429), .b(gnd), .g(inst[13]));
NEMR4T g283(.s(AA_429), .d(AA_442), .b(vdd), .g(irq));
NEMR4T g284(.s(AA_429), .d(AA_393), .b(gnd), .g(irq));
NEMR4T g285(.s(AA_182), .d(AA_180), .b(gnd), .g(inst[16]));
NEMR4T g286(.s(AA_180), .d(AA_171), .b(vdd), .g(inst[13]));
NEMR4T g287(.s(AA_171), .d(AA_170), .b(vdd), .g(irq));
NEMR4T g288(.s(AA_170), .d(AA_430), .b(gnd), .g(inst[17]));
NEMR4T g289(.s(AA_430), .d(AA_397), .b(vdd), .g(ireset));
NEMR4T g290(.s(AA_171), .d(AA_150), .b(gnd), .g(irq));
NEMR4T g291(.s(AA_150), .d(AA_393), .b(vdd), .g(inst[17]));
NEMR4T g292(.s(AA_150), .d(AA_111), .b(gnd), .g(inst[17]));
NEMR4T g293(.s(AA_111), .d(AA_393), .b(vdd), .g(ireset));
NEMR4T g294(.s(AA_111), .d(AA_391), .b(gnd), .g(ireset));
NEMR4T g295(.s(BB_100_30), .d(AA_431), .b(vdd), .g(inst[16]));
NEMR4T g296(.s(AA_431), .d(AA_429), .b(vdd), .g(inst[13]));
NEMR4T g297(.s(BB_100_30), .d(BB_100_30222221), .b(gnd), .g(inst[16]));
NEMR4T g298(.s(BB_100_30222221), .d(AA_169), .b(vdd), .g(inst[13]));
NEMR4T g299(.s(BB_100_30222221), .d(AA_153), .b(gnd), .g(inst[13]));
NEMR4T g300(.s(AA_153), .d(AA_117), .b(vdd), .g(irq));
NEMR4T g301(.s(AA_117), .d(AA_430), .b(gnd), .g(inst[17]));
NEMR4T g302(.s(AA_117), .d(AA_393), .b(gnd), .g(ireset));
NEMR4T g303(.s(AA_153), .d(AA_150), .b(gnd), .g(irq));
NEMR4T g304(.s(pcsel[1]), .d(BB_100_31), .b(gnd), .g(inst[12]));
NEMR4T g305(.s(BB_100_31), .d(BB_100_310), .b(vdd), .g(z));
NEMR4T g306(.s(BB_100_310), .d(AA_181), .b(vdd), .g(c));
NEMR4T g307(.s(AA_181), .d(AA_173), .b(vdd), .g(inst[10]));
NEMR4T g308(.s(AA_173), .d(AA_154), .b(vdd), .g(inst[14]));
NEMR4T g309(.s(AA_154), .d(AA_169), .b(gnd), .g(inst[16]));
NEMR4T g310(.s(AA_173), .d(AA_462), .b(gnd), .g(inst[14]));
NEMR4T g311(.s(AA_462), .d(AA_455), .b(gnd), .g(inst[16]));
NEMR4T g312(.s(AA_455), .d(AA_432), .b(vdd), .g(inst[13]));
NEMR4T g313(.s(AA_432), .d(AA_401), .b(vdd), .g(irq));
NEMR4T g314(.s(AA_432), .d(AA_393), .b(gnd), .g(irq));
NEMR4T g315(.s(AA_173), .d(AA_429), .b(vdd), .g(inst[16]));
NEMR4T g316(.s(AA_181), .d(AA_176), .b(gnd), .g(inst[10]));
NEMR4T g317(.s(AA_176), .d(AA_179), .b(vdd), .g(inst[14]));
NEMR4T g318(.s(AA_176), .d(AA_431), .b(vdd), .g(inst[16]));
NEMR4T g319(.s(AA_176), .d(AA_125), .b(gnd), .g(inst[16]));
NEMR4T g320(.s(AA_125), .d(AA_169), .b(vdd), .g(inst[13]));
NEMR4T g321(.s(BB_100_310), .d(BB_100_3101), .b(gnd), .g(c));
NEMR4T g322(.s(BB_100_3101), .d(AA_181), .b(vdd), .g(inst[11]));
NEMR4T g323(.s(BB_100_3101), .d(BB_100_31011), .b(gnd), .g(inst[11]));
NEMR4T g324(.s(BB_100_31011), .d(AA_162), .b(gnd), .g(inst[10]));
NEMR4T g325(.s(AA_162), .d(AA_129), .b(vdd), .g(inst[14]));
NEMR4T g326(.s(AA_129), .d(AA_429), .b(vdd), .g(inst[16]));
NEMR4T g327(.s(AA_129), .d(AA_169), .b(gnd), .g(inst[16]));
NEMR4T g328(.s(BB_100_310), .d(BB_100_310221), .b(gnd), .g(inst[10]));
NEMR4T g329(.s(BB_100_310221), .d(AA_182), .b(gnd), .g(inst[14]));
NEMR4T g330(.s(BB_100_310), .d(AA_164), .b(gnd), .g(inst[16]));
NEMR4T g331(.s(AA_164), .d(AA_153), .b(gnd), .g(inst[13]));
NEMR4T g332(.s(BB_100_31), .d(BB_100_311), .b(gnd), .g(z));
NEMR4T g333(.s(BB_100_311), .d(BB_100_3110), .b(vdd), .g(c));
NEMR4T g334(.s(BB_100_3110), .d(BB_100_31101), .b(gnd), .g(inst[11]));
NEMR4T g335(.s(BB_100_31101), .d(AA_173), .b(vdd), .g(inst[10]));
NEMR4T g336(.s(BB_100_31101), .d(BB_100_311011), .b(gnd), .g(inst[10]));
NEMR4T g337(.s(BB_100_311011), .d(AA_179), .b(vdd), .g(inst[14]));
NEMR4T g338(.s(BB_100_3110), .d(AA_165), .b(gnd), .g(inst[10]));
NEMR4T g339(.s(AA_165), .d(AA_136), .b(gnd), .g(inst[14]));
NEMR4T g340(.s(AA_136), .d(AA_431), .b(vdd), .g(inst[16]));
NEMR4T g341(.s(AA_136), .d(AA_125), .b(gnd), .g(inst[16]));
NEMR4T g342(.s(BB_100_3110), .d(AA_164), .b(gnd), .g(inst[16]));
NEMR4T g343(.s(BB_100_311), .d(BB_100_3111), .b(gnd), .g(c));
NEMR4T g344(.s(BB_100_3111), .d(BB_100_31110), .b(vdd), .g(inst[11]));
NEMR4T g345(.s(BB_100_31110), .d(AA_165), .b(gnd), .g(inst[10]));
NEMR4T g346(.s(BB_100_31110), .d(AA_164), .b(gnd), .g(inst[16]));
NEMR4T g347(.s(BB_100_3111), .d(BB_100_31111), .b(gnd), .g(inst[11]));
NEMR4T g348(.s(BB_100_31111), .d(AA_139), .b(vdd), .g(inst[10]));
NEMR4T g349(.s(AA_139), .d(AA_164), .b(gnd), .g(inst[16]));
NEMR4T g350(.s(BB_100_31111), .d(BB_100_311111), .b(gnd), .g(inst[10]));
NEMR4T g351(.s(BB_100_311111), .d(AA_148), .b(vdd), .g(inst[14]));
NEMR4T g352(.s(BB_100_311111), .d(AA_139), .b(gnd), .g(inst[14]));
NEMR4T g353(.s(BB_100_311), .d(BB_100_31120), .b(vdd), .g(inst[11]));
NEMR4T g354(.s(BB_100_31120), .d(AA_176), .b(vdd), .g(inst[10]));
NEMR4T g355(.s(BB_100_31120), .d(AA_162), .b(gnd), .g(inst[10]));
NEMR4T g356(.s(BB_100_31120), .d(AA_182), .b(gnd), .g(inst[14]));
NEMR4T g357(.s(BB_100_311), .d(BB_100_31121), .b(gnd), .g(inst[11]));
NEMR4T g358(.s(BB_100_31121), .d(BB_100_311211), .b(gnd), .g(inst[10]));
NEMR4T g359(.s(BB_100_311211), .d(AA_136), .b(vdd), .g(inst[14]));
NEMR4T g360(.s(BB_100_311211), .d(AA_182), .b(gnd), .g(inst[14]));
NEMR4T g361(.s(BB_100_31), .d(BB_100_3121), .b(gnd), .g(c));
NEMR4T g362(.s(BB_100_3121), .d(BB_100_31211), .b(gnd), .g(inst[11]));
NEMR4T g363(.s(BB_100_31211), .d(BB_100_312110), .b(vdd), .g(inst[10]));
NEMR4T g364(.s(BB_100_312110), .d(AA_179), .b(vdd), .g(inst[14]));
NEMR4T g365(.s(BB_100_312110), .d(AA_182), .b(gnd), .g(inst[14]));
NEMR4T g366(.s(BB_100_312110), .d(AA_431), .b(vdd), .g(inst[16]));
NEMR4T g367(.s(BB_100_312110), .d(AA_125), .b(gnd), .g(inst[16]));
NEMR4T g368(.s(BB_100_31211), .d(AA_165), .b(gnd), .g(inst[10]));
NEMR4T g369(.s(pcsel[1]), .d(BB_100_3222220), .b(vdd), .g(inst[14]));
NEMR4T g370(.s(BB_100_3222220), .d(BB_100_32222201), .b(gnd), .g(inst[16]));
NEMR4T g371(.s(BB_100_32222201), .d(AA_167), .b(vdd), .g(inst[13]));
NEMR4T g372(.s(pcsel[1]), .d(BB_100_3222221), .b(gnd), .g(inst[14]));
NEMR4T g373(.s(BB_100_3222221), .d(BB_100_32222211), .b(gnd), .g(inst[16]));
NEMR4T g374(.s(BB_100_32222211), .d(AA_433), .b(vdd), .g(inst[13]));
NEMR4T g375(.s(AA_433), .d(AA_425), .b(vdd), .g(irq));
NEMR4T g376(.s(BB_100_32222211), .d(AA_169), .b(gnd), .g(inst[13]));
NEMR4T g377(.s(pcsel[0]), .d(AA_231), .b(vdd), .g(inst[12]));
NEMR4T g378(.s(AA_231), .d(AA_429), .b(vdd), .g(inst[16]));
NEMR4T g379(.s(AA_231), .d(AA_227), .b(gnd), .g(inst[16]));
NEMR4T g380(.s(AA_227), .d(AA_224), .b(vdd), .g(inst[13]));
NEMR4T g381(.s(AA_224), .d(AA_441), .b(vdd), .g(irq));
NEMR4T g382(.s(AA_224), .d(AA_424), .b(gnd), .g(irq));
NEMR4T g383(.s(AA_224), .d(AA_425), .b(vdd), .g(inst[17]));
NEMR4T g384(.s(AA_224), .d(AA_428), .b(gnd), .g(inst[17]));
NEMR4T g385(.s(AA_227), .d(AA_225), .b(gnd), .g(inst[13]));
NEMR4T g386(.s(AA_225), .d(AA_214), .b(vdd), .g(irq));
NEMR4T g387(.s(AA_214), .d(AA_427), .b(gnd), .g(inst[17]));
NEMR4T g388(.s(AA_214), .d(AA_393), .b(gnd), .g(ireset));
NEMR4T g389(.s(AA_225), .d(AA_215), .b(gnd), .g(irq));
NEMR4T g390(.s(AA_215), .d(AA_393), .b(vdd), .g(inst[17]));
NEMR4T g391(.s(AA_215), .d(AA_191), .b(gnd), .g(inst[17]));
NEMR4T g392(.s(AA_191), .d(AA_393), .b(vdd), .g(ireset));
NEMR4T g393(.s(AA_191), .d(AA_394), .b(gnd), .g(ireset));
NEMR4T g394(.s(AA_227), .d(AA_226), .b(vdd), .g(irq));
NEMR4T g395(.s(AA_226), .d(AA_401), .b(vdd), .g(inst[17]));
NEMR4T g396(.s(AA_226), .d(AA_430), .b(gnd), .g(inst[17]));
NEMR4T g397(.s(AA_227), .d(AA_217), .b(gnd), .g(irq));
NEMR4T g398(.s(AA_217), .d(AA_426), .b(gnd), .g(inst[17]));
NEMR4T g399(.s(pcsel[0]), .d(BB_183_31), .b(gnd), .g(inst[12]));
NEMR4T g400(.s(BB_183_31), .d(BB_183_310), .b(vdd), .g(z));
NEMR4T g401(.s(BB_183_310), .d(AA_232), .b(vdd), .g(c));
NEMR4T g402(.s(AA_232), .d(AA_429), .b(vdd), .g(inst[10]));
NEMR4T g403(.s(AA_232), .d(AA_228), .b(gnd), .g(inst[10]));
NEMR4T g404(.s(AA_228), .d(AA_220), .b(gnd), .g(inst[16]));
NEMR4T g405(.s(AA_220), .d(AA_224), .b(vdd), .g(inst[13]));
NEMR4T g406(.s(AA_220), .d(AA_226), .b(vdd), .g(irq));
NEMR4T g407(.s(AA_220), .d(AA_217), .b(gnd), .g(irq));
NEMR4T g408(.s(BB_183_310), .d(BB_183_3101), .b(gnd), .g(c));
NEMR4T g409(.s(BB_183_3101), .d(AA_232), .b(vdd), .g(inst[11]));
NEMR4T g410(.s(BB_183_3101), .d(BB_183_31011), .b(gnd), .g(inst[11]));
NEMR4T g411(.s(BB_183_31011), .d(AA_462), .b(gnd), .g(inst[10]));
NEMR4T g412(.s(BB_183_310), .d(BB_183_310221), .b(gnd), .g(inst[10]));
NEMR4T g413(.s(BB_183_310221), .d(AA_429), .b(vdd), .g(inst[16]));
NEMR4T g414(.s(BB_183_310221), .d(AA_229), .b(gnd), .g(inst[16]));
NEMR4T g415(.s(AA_229), .d(AA_225), .b(gnd), .g(inst[13]));
NEMR4T g416(.s(BB_183_31), .d(BB_183_311), .b(gnd), .g(z));
NEMR4T g417(.s(BB_183_311), .d(BB_183_3110), .b(vdd), .g(c));
NEMR4T g418(.s(BB_183_3110), .d(BB_183_31101), .b(gnd), .g(inst[11]));
NEMR4T g419(.s(BB_183_31101), .d(AA_429), .b(vdd), .g(inst[10]));
NEMR4T g420(.s(BB_183_31101), .d(BB_183_311011), .b(gnd), .g(inst[10]));
NEMR4T g421(.s(BB_183_311011), .d(BB_183_3110111), .b(gnd), .g(inst[16]));
NEMR4T g422(.s(BB_183_3110111), .d(AA_224), .b(vdd), .g(inst[13]));
NEMR4T g423(.s(BB_183_3110), .d(AA_230), .b(gnd), .g(inst[10]));
NEMR4T g424(.s(AA_230), .d(AA_223), .b(gnd), .g(inst[16]));
NEMR4T g425(.s(AA_223), .d(AA_207), .b(gnd), .g(inst[13]));
NEMR4T g426(.s(AA_207), .d(AA_226), .b(vdd), .g(irq));
NEMR4T g427(.s(AA_207), .d(AA_217), .b(gnd), .g(irq));
NEMR4T g428(.s(BB_183_311), .d(BB_183_3111), .b(gnd), .g(c));
NEMR4T g429(.s(BB_183_3111), .d(BB_183_31110), .b(vdd), .g(inst[11]));
NEMR4T g430(.s(BB_183_31110), .d(AA_230), .b(gnd), .g(inst[10]));
NEMR4T g431(.s(BB_183_3111), .d(BB_183_31111), .b(gnd), .g(inst[11]));
NEMR4T g432(.s(BB_183_31111), .d(BB_183_311111), .b(gnd), .g(inst[10]));
NEMR4T g433(.s(BB_183_311111), .d(BB_183_3111111), .b(gnd), .g(inst[16]));
NEMR4T g434(.s(BB_183_3111111), .d(BB_183_31111110), .b(vdd), .g(inst[13]));
NEMR4T g435(.s(BB_183_31111110), .d(BB_183_311111100), .b(vdd), .g(irq));
NEMR4T g436(.s(BB_183_311111100), .d(AA_427), .b(gnd), .g(inst[17]));
NEMR4T g437(.s(BB_183_31111110), .d(AA_215), .b(gnd), .g(irq));
NEMR4T g438(.s(BB_183_311), .d(BB_183_31120), .b(vdd), .g(inst[11]));
NEMR4T g439(.s(BB_183_31120), .d(AA_228), .b(vdd), .g(inst[10]));
NEMR4T g440(.s(BB_183_31120), .d(BB_183_311201), .b(gnd), .g(inst[10]));
NEMR4T g441(.s(BB_183_311201), .d(AA_431), .b(gnd), .g(inst[16]));
NEMR4T g442(.s(BB_183_31120), .d(AA_429), .b(vdd), .g(inst[16]));
NEMR4T g443(.s(BB_183_31120), .d(AA_229), .b(gnd), .g(inst[16]));
NEMR4T g444(.s(BB_183_311), .d(BB_183_31121), .b(gnd), .g(inst[11]));
NEMR4T g445(.s(BB_183_31121), .d(BB_183_311211), .b(gnd), .g(inst[10]));
NEMR4T g446(.s(BB_183_311211), .d(AA_429), .b(vdd), .g(inst[16]));
NEMR4T g447(.s(BB_183_311211), .d(BB_183_3112111), .b(gnd), .g(inst[16]));
NEMR4T g448(.s(BB_183_3112111), .d(AA_207), .b(vdd), .g(inst[13]));
NEMR4T g449(.s(BB_183_3112111), .d(AA_225), .b(gnd), .g(inst[13]));
NEMR4T g450(.s(BB_183_31), .d(BB_183_3121), .b(gnd), .g(c));
NEMR4T g451(.s(BB_183_3121), .d(BB_183_31211), .b(gnd), .g(inst[11]));
NEMR4T g452(.s(BB_183_31211), .d(AA_231), .b(vdd), .g(inst[10]));
NEMR4T g453(.s(BB_183_31211), .d(BB_183_312111), .b(gnd), .g(inst[10]));
NEMR4T g454(.s(BB_183_312111), .d(BB_183_3121111), .b(gnd), .g(inst[16]));
NEMR4T g455(.s(BB_183_3121111), .d(AA_433), .b(vdd), .g(inst[13]));
NEMR4T g456(.s(BB_183_3121111), .d(AA_207), .b(gnd), .g(inst[13]));
NEMR4T g457(.s(stsel[0]), .d(AA_284), .b(vdd), .g(inst[12]));
NEMR4T g458(.s(AA_284), .d(AA_280), .b(vdd), .g(inst[14]));
NEMR4T g459(.s(AA_280), .d(AA_273), .b(gnd), .g(inst[16]));
NEMR4T g460(.s(AA_273), .d(AA_272), .b(vdd), .g(inst[13]));
NEMR4T g461(.s(AA_272), .d(AA_434), .b(vdd), .g(irq));
NEMR4T g462(.s(AA_434), .d(AA_397), .b(gnd), .g(inst[17]));
NEMR4T g463(.s(AA_272), .d(AA_260), .b(gnd), .g(inst[17]));
NEMR4T g464(.s(AA_260), .d(AA_391), .b(vdd), .g(ireset));
NEMR4T g465(.s(AA_260), .d(AA_395), .b(gnd), .g(ireset));
NEMR4T g466(.s(AA_273), .d(AA_404), .b(vdd), .g(irq));
NEMR4T g467(.s(AA_273), .d(AA_262), .b(gnd), .g(irq));
NEMR4T g468(.s(AA_262), .d(AA_435), .b(vdd), .g(inst[17]));
NEMR4T g469(.s(AA_435), .d(AA_393), .b(vdd), .g(ireset));
NEMR4T g470(.s(AA_435), .d(AA_392), .b(gnd), .g(ireset));
NEMR4T g471(.s(AA_262), .d(AA_241), .b(gnd), .g(inst[17]));
NEMR4T g472(.s(AA_241), .d(AA_394), .b(vdd), .g(ireset));
NEMR4T g473(.s(AA_241), .d(AA_397), .b(gnd), .g(ireset));
NEMR4T g474(.s(AA_284), .d(AA_281), .b(gnd), .g(inst[14]));
NEMR4T g475(.s(AA_281), .d(AA_274), .b(gnd), .g(inst[16]));
NEMR4T g476(.s(AA_274), .d(AA_242), .b(vdd), .g(inst[13]));
NEMR4T g477(.s(AA_242), .d(AA_392), .b(vdd), .g(irq));
NEMR4T g478(.s(AA_242), .d(AA_435), .b(gnd), .g(irq));
NEMR4T g479(.s(AA_274), .d(AA_263), .b(gnd), .g(inst[13]));
NEMR4T g480(.s(AA_263), .d(AA_404), .b(vdd), .g(irq));
NEMR4T g481(.s(AA_263), .d(AA_262), .b(gnd), .g(irq));
NEMR4T g482(.s(AA_284), .d(AA_242), .b(vdd), .g(inst[16]));
NEMR4T g483(.s(AA_284), .d(AA_282), .b(gnd), .g(inst[16]));
NEMR4T g484(.s(AA_282), .d(AA_275), .b(gnd), .g(inst[13]));
NEMR4T g485(.s(AA_275), .d(AA_245), .b(vdd), .g(irq));
NEMR4T g486(.s(AA_245), .d(AA_392), .b(gnd), .g(inst[17]));
NEMR4T g487(.s(AA_275), .d(AA_264), .b(gnd), .g(irq));
NEMR4T g488(.s(AA_264), .d(AA_260), .b(gnd), .g(inst[17]));
NEMR4T g489(.s(stsel[0]), .d(BB_233_31), .b(gnd), .g(inst[12]));
NEMR4T g490(.s(BB_233_31), .d(BB_233_310), .b(vdd), .g(z));
NEMR4T g491(.s(BB_233_310), .d(AA_285), .b(vdd), .g(c));
NEMR4T g492(.s(AA_285), .d(AA_242), .b(vdd), .g(inst[10]));
NEMR4T g493(.s(AA_285), .d(AA_283), .b(gnd), .g(inst[10]));
NEMR4T g494(.s(AA_283), .d(AA_280), .b(vdd), .g(inst[14]));
NEMR4T g495(.s(AA_283), .d(AA_242), .b(vdd), .g(inst[16]));
NEMR4T g496(.s(AA_283), .d(AA_282), .b(gnd), .g(inst[16]));
NEMR4T g497(.s(BB_233_310), .d(BB_233_3101), .b(gnd), .g(c));
NEMR4T g498(.s(BB_233_3101), .d(AA_285), .b(vdd), .g(inst[11]));
NEMR4T g499(.s(BB_233_3101), .d(BB_233_31011), .b(gnd), .g(inst[11]));
NEMR4T g500(.s(BB_233_31011), .d(AA_253), .b(gnd), .g(inst[10]));
NEMR4T g501(.s(AA_253), .d(AA_242), .b(vdd), .g(inst[14]));
NEMR4T g502(.s(BB_233_310), .d(BB_233_310221), .b(gnd), .g(inst[10]));
NEMR4T g503(.s(BB_233_310221), .d(AA_281), .b(gnd), .g(inst[14]));
NEMR4T g504(.s(BB_233_31), .d(BB_233_311), .b(gnd), .g(z));
NEMR4T g505(.s(BB_233_311), .d(BB_233_3110), .b(vdd), .g(c));
NEMR4T g506(.s(BB_233_3110), .d(BB_233_31101), .b(gnd), .g(inst[11]));
NEMR4T g507(.s(BB_233_31101), .d(AA_242), .b(vdd), .g(inst[10]));
NEMR4T g508(.s(BB_233_31101), .d(BB_233_311011), .b(gnd), .g(inst[10]));
NEMR4T g509(.s(BB_233_311011), .d(AA_280), .b(vdd), .g(inst[14]));
NEMR4T g510(.s(BB_233_3110), .d(AA_279), .b(gnd), .g(inst[10]));
NEMR4T g511(.s(AA_279), .d(AA_269), .b(gnd), .g(inst[14]));
NEMR4T g512(.s(AA_269), .d(AA_242), .b(vdd), .g(inst[16]));
NEMR4T g513(.s(AA_269), .d(AA_282), .b(gnd), .g(inst[16]));
NEMR4T g514(.s(BB_233_311), .d(BB_233_3111), .b(gnd), .g(c));
NEMR4T g515(.s(BB_233_3111), .d(BB_233_31110), .b(vdd), .g(inst[11]));
NEMR4T g516(.s(BB_233_31110), .d(AA_279), .b(gnd), .g(inst[10]));
NEMR4T g517(.s(BB_233_3111), .d(BB_233_31111), .b(gnd), .g(inst[11]));
NEMR4T g518(.s(BB_233_31111), .d(BB_233_311111), .b(gnd), .g(inst[10]));
NEMR4T g519(.s(BB_233_311111), .d(AA_281), .b(vdd), .g(inst[14]));
NEMR4T g520(.s(BB_233_311), .d(BB_233_31120), .b(vdd), .g(inst[11]));
NEMR4T g521(.s(BB_233_31120), .d(AA_283), .b(vdd), .g(inst[10]));
NEMR4T g522(.s(BB_233_31120), .d(AA_253), .b(gnd), .g(inst[10]));
NEMR4T g523(.s(BB_233_31120), .d(AA_281), .b(gnd), .g(inst[14]));
NEMR4T g524(.s(BB_233_311), .d(BB_233_31121), .b(gnd), .g(inst[11]));
NEMR4T g525(.s(BB_233_31121), .d(BB_233_311211), .b(gnd), .g(inst[10]));
NEMR4T g526(.s(BB_233_311211), .d(AA_269), .b(vdd), .g(inst[14]));
NEMR4T g527(.s(BB_233_311211), .d(AA_281), .b(gnd), .g(inst[14]));
NEMR4T g528(.s(BB_233_31), .d(BB_233_3121), .b(gnd), .g(c));
NEMR4T g529(.s(BB_233_3121), .d(BB_233_31211), .b(gnd), .g(inst[11]));
NEMR4T g530(.s(BB_233_31211), .d(AA_284), .b(vdd), .g(inst[10]));
NEMR4T g531(.s(BB_233_31211), .d(AA_279), .b(gnd), .g(inst[10]));
NEMR4T g532(.s(stsel[1]), .d(BB_286_30), .b(vdd), .g(inst[12]));
NEMR4T g533(.s(BB_286_30), .d(AA_341), .b(vdd), .g(inst[14]));
NEMR4T g534(.s(AA_341), .d(AA_456), .b(vdd), .g(inst[16]));
NEMR4T g535(.s(AA_456), .d(AA_436), .b(gnd), .g(inst[13]));
NEMR4T g536(.s(AA_436), .d(AA_419), .b(vdd), .g(irq));
NEMR4T g537(.s(AA_436), .d(AA_392), .b(vdd), .g(inst[17]));
NEMR4T g538(.s(AA_436), .d(AA_403), .b(gnd), .g(inst[17]));
NEMR4T g539(.s(AA_341), .d(AA_461), .b(gnd), .g(inst[13]));
NEMR4T g540(.s(BB_286_30), .d(AA_342), .b(gnd), .g(inst[14]));
NEMR4T g541(.s(AA_342), .d(AA_292), .b(vdd), .g(inst[16]));
NEMR4T g542(.s(AA_292), .d(AA_392), .b(gnd), .g(inst[13]));
NEMR4T g543(.s(AA_342), .d(AA_340), .b(gnd), .g(inst[16]));
NEMR4T g544(.s(AA_340), .d(AA_451), .b(vdd), .g(inst[13]));
NEMR4T g545(.s(BB_286_30), .d(AA_294), .b(vdd), .g(inst[16]));
NEMR4T g546(.s(AA_294), .d(AA_392), .b(vdd), .g(inst[13]));
NEMR4T g547(.s(BB_286_30), .d(BB_286_30222221), .b(gnd), .g(inst[16]));
NEMR4T g548(.s(BB_286_30222221), .d(AA_461), .b(vdd), .g(inst[13]));
NEMR4T g549(.s(BB_286_30222221), .d(AA_451), .b(gnd), .g(inst[13]));
NEMR4T g550(.s(stsel[1]), .d(BB_286_31), .b(gnd), .g(inst[12]));
NEMR4T g551(.s(BB_286_31), .d(BB_286_310), .b(vdd), .g(z));
NEMR4T g552(.s(BB_286_310), .d(AA_336), .b(vdd), .g(c));
NEMR4T g553(.s(AA_336), .d(AA_335), .b(vdd), .g(inst[10]));
NEMR4T g554(.s(AA_335), .d(AA_334), .b(vdd), .g(inst[14]));
NEMR4T g555(.s(AA_334), .d(AA_461), .b(gnd), .g(inst[16]));
NEMR4T g556(.s(AA_335), .d(AA_298), .b(gnd), .g(inst[14]));
NEMR4T g557(.s(AA_298), .d(AA_294), .b(gnd), .g(inst[16]));
NEMR4T g558(.s(AA_335), .d(AA_392), .b(vdd), .g(inst[16]));
NEMR4T g559(.s(AA_336), .d(AA_325), .b(gnd), .g(inst[10]));
NEMR4T g560(.s(AA_325), .d(AA_341), .b(vdd), .g(inst[14]));
NEMR4T g561(.s(AA_325), .d(AA_294), .b(vdd), .g(inst[16]));
NEMR4T g562(.s(AA_325), .d(AA_302), .b(gnd), .g(inst[16]));
NEMR4T g563(.s(AA_302), .d(AA_461), .b(vdd), .g(inst[13]));
NEMR4T g564(.s(BB_286_310), .d(BB_286_3101), .b(gnd), .g(c));
NEMR4T g565(.s(BB_286_3101), .d(AA_336), .b(vdd), .g(inst[11]));
NEMR4T g566(.s(BB_286_3101), .d(BB_286_31011), .b(gnd), .g(inst[11]));
NEMR4T g567(.s(BB_286_31011), .d(AA_326), .b(gnd), .g(inst[10]));
NEMR4T g568(.s(AA_326), .d(AA_308), .b(vdd), .g(inst[14]));
NEMR4T g569(.s(AA_308), .d(AA_392), .b(vdd), .g(inst[16]));
NEMR4T g570(.s(AA_308), .d(AA_461), .b(gnd), .g(inst[16]));
NEMR4T g571(.s(BB_286_310), .d(BB_286_310221), .b(gnd), .g(inst[10]));
NEMR4T g572(.s(BB_286_310221), .d(AA_342), .b(gnd), .g(inst[14]));
NEMR4T g573(.s(BB_286_310), .d(AA_460), .b(gnd), .g(inst[16]));
NEMR4T g574(.s(BB_286_31), .d(BB_286_311), .b(gnd), .g(z));
NEMR4T g575(.s(BB_286_311), .d(BB_286_3110), .b(vdd), .g(c));
NEMR4T g576(.s(BB_286_3110), .d(BB_286_31101), .b(gnd), .g(inst[11]));
NEMR4T g577(.s(BB_286_31101), .d(AA_335), .b(vdd), .g(inst[10]));
NEMR4T g578(.s(BB_286_31101), .d(BB_286_311011), .b(gnd), .g(inst[10]));
NEMR4T g579(.s(BB_286_311011), .d(AA_341), .b(vdd), .g(inst[14]));
NEMR4T g580(.s(BB_286_3110), .d(AA_328), .b(gnd), .g(inst[10]));
NEMR4T g581(.s(AA_328), .d(AA_311), .b(gnd), .g(inst[14]));
NEMR4T g582(.s(AA_311), .d(AA_294), .b(vdd), .g(inst[16]));
NEMR4T g583(.s(AA_311), .d(AA_302), .b(gnd), .g(inst[16]));
NEMR4T g584(.s(BB_286_3110), .d(AA_460), .b(gnd), .g(inst[16]));
NEMR4T g585(.s(BB_286_311), .d(BB_286_3111), .b(gnd), .g(c));
NEMR4T g586(.s(BB_286_3111), .d(BB_286_31110), .b(vdd), .g(inst[11]));
NEMR4T g587(.s(BB_286_31110), .d(AA_328), .b(gnd), .g(inst[10]));
NEMR4T g588(.s(BB_286_31110), .d(AA_460), .b(gnd), .g(inst[16]));
NEMR4T g589(.s(BB_286_3111), .d(BB_286_31111), .b(gnd), .g(inst[11]));
NEMR4T g590(.s(BB_286_31111), .d(AA_313), .b(vdd), .g(inst[10]));
NEMR4T g591(.s(AA_313), .d(AA_460), .b(gnd), .g(inst[16]));
NEMR4T g592(.s(BB_286_31111), .d(BB_286_311111), .b(gnd), .g(inst[10]));
NEMR4T g593(.s(BB_286_311111), .d(AA_292), .b(vdd), .g(inst[14]));
NEMR4T g594(.s(BB_286_311111), .d(AA_313), .b(gnd), .g(inst[14]));
NEMR4T g595(.s(BB_286_311), .d(BB_286_31120), .b(vdd), .g(inst[11]));
NEMR4T g596(.s(BB_286_31120), .d(AA_325), .b(vdd), .g(inst[10]));
NEMR4T g597(.s(BB_286_31120), .d(AA_326), .b(gnd), .g(inst[10]));
NEMR4T g598(.s(BB_286_31120), .d(AA_342), .b(gnd), .g(inst[14]));
NEMR4T g599(.s(BB_286_311), .d(BB_286_31121), .b(gnd), .g(inst[11]));
NEMR4T g600(.s(BB_286_31121), .d(BB_286_311211), .b(gnd), .g(inst[10]));
NEMR4T g601(.s(BB_286_311211), .d(AA_311), .b(vdd), .g(inst[14]));
NEMR4T g602(.s(BB_286_311211), .d(AA_342), .b(gnd), .g(inst[14]));
NEMR4T g603(.s(BB_286_31), .d(BB_286_3121), .b(gnd), .g(c));
NEMR4T g604(.s(BB_286_3121), .d(BB_286_31211), .b(gnd), .g(inst[11]));
NEMR4T g605(.s(BB_286_31211), .d(BB_286_312110), .b(vdd), .g(inst[10]));
NEMR4T g606(.s(BB_286_312110), .d(AA_341), .b(vdd), .g(inst[14]));
NEMR4T g607(.s(BB_286_312110), .d(AA_342), .b(gnd), .g(inst[14]));
NEMR4T g608(.s(BB_286_312110), .d(AA_294), .b(vdd), .g(inst[16]));
NEMR4T g609(.s(BB_286_312110), .d(AA_302), .b(gnd), .g(inst[16]));
NEMR4T g610(.s(BB_286_31211), .d(AA_328), .b(gnd), .g(inst[10]));
NEMR4T g611(.s(stsel[1]), .d(BB_286_3222220), .b(vdd), .g(inst[14]));
NEMR4T g612(.s(BB_286_3222220), .d(BB_286_32222201), .b(gnd), .g(inst[16]));
NEMR4T g613(.s(BB_286_32222201), .d(AA_436), .b(vdd), .g(inst[13]));
NEMR4T g614(.s(stsel[1]), .d(BB_286_3222221), .b(gnd), .g(inst[14]));
NEMR4T g615(.s(BB_286_3222221), .d(BB_286_32222211), .b(gnd), .g(inst[16]));
NEMR4T g616(.s(BB_286_32222211), .d(AA_461), .b(gnd), .g(inst[13]));
NEMR4T g617(.s(read_strobe), .d(AA_392), .b(vdd), .g(inst[14]));
NEMR4T g618(.s(read_strobe), .d(BB_343_31), .b(gnd), .g(inst[14]));
NEMR4T g619(.s(BB_343_31), .d(BB_343_310), .b(vdd), .g(inst[16]));
NEMR4T g620(.s(BB_343_310), .d(BB_343_3100), .b(vdd), .g(inst[13]));
NEMR4T g621(.s(BB_343_3100), .d(AA_402), .b(vdd), .g(irq));
NEMR4T g622(.s(BB_343_3100), .d(AA_423), .b(gnd), .g(inst[17]));
NEMR4T g623(.s(BB_343_310), .d(AA_420), .b(gnd), .g(irq));
NEMR4T g624(.s(BB_343_31), .d(BB_343_311), .b(gnd), .g(inst[16]));
NEMR4T g625(.s(BB_343_311), .d(AA_392), .b(vdd), .g(inst[13]));
NEMR4T g626(.s(BB_343_311), .d(AA_453), .b(gnd), .g(inst[13]));
NEMR4T g627(.s(BB_343_31), .d(BB_343_3121), .b(gnd), .g(inst[13]));
NEMR4T g628(.s(BB_343_3121), .d(AA_392), .b(vdd), .g(irq));
NEMR4T g629(.s(BB_343_3121), .d(BB_343_31211), .b(gnd), .g(irq));
NEMR4T g630(.s(BB_343_31211), .d(AA_423), .b(gnd), .g(inst[17]));
NEMR4T g631(.s(write_strobe), .d(BB_350_30), .b(vdd), .g(clk));
NEMR4T g632(.s(BB_350_30), .d(BB_350_301), .b(gnd), .g(inst[14]));
NEMR4T g633(.s(BB_350_301), .d(BB_350_3010), .b(vdd), .g(inst[16]));
NEMR4T g634(.s(BB_350_3010), .d(AA_436), .b(vdd), .g(inst[13]));
NEMR4T g635(.s(BB_350_3010), .d(AA_452), .b(gnd), .g(irq));
NEMR4T g636(.s(BB_350_301), .d(AA_451), .b(gnd), .g(inst[13]));
NEMR4T g637(.s(write_strobe), .d(BB_350_31), .b(gnd), .g(clk));
NEMR4T g638(.s(BB_350_31), .d(BB_350_311), .b(gnd), .g(inst[14]));
NEMR4T g639(.s(BB_350_311), .d(AA_392), .b(vdd), .g(inst[16]));
NEMR4T g640(.s(BB_350_311), .d(AA_460), .b(gnd), .g(inst[16]));
NEMR4T g641(.s(write_strobe), .d(AA_392), .b(vdd), .g(inst[14]));
NEMR4T g642(.s(write_strobe), .d(BB_350_321), .b(gnd), .g(inst[14]));
NEMR4T g643(.s(BB_350_321), .d(AA_464), .b(gnd), .g(inst[16]));
NEMR4T g644(.s(interrupt_ack), .d(AA_392), .b(vdd), .g(irq));
NEMR4T g645(.s(interrupt_ack), .d(BB_360_31), .b(gnd), .g(irq));
NEMR4T g646(.s(BB_360_31), .d(vdd), .b(vdd), .g(ireset));
NEMR4T g647(.s(BB_360_31), .d(gnd), .b(gnd), .g(ireset));
NEMR4T g648(.s(next_interrupt_enabled), .d(BB_361_30), .b(vdd), .g(interrupt_enabled));
NEMR4T g649(.s(BB_361_30), .d(AA_392), .b(vdd), .g(inst[0]));
NEMR4T g650(.s(BB_361_30), .d(BB_361_301), .b(gnd), .g(inst[0]));
NEMR4T g651(.s(BB_361_301), .d(AA_392), .b(vdd), .g(inst[16]));
NEMR4T g652(.s(BB_361_301), .d(BB_361_3011), .b(gnd), .g(inst[16]));
NEMR4T g653(.s(BB_361_3011), .d(BB_361_30110), .b(vdd), .g(inst[13]));
NEMR4T g654(.s(BB_361_30110), .d(BB_361_301100), .b(vdd), .g(irq));
NEMR4T g655(.s(BB_361_301100), .d(AA_395), .b(gnd), .g(inst[17]));
NEMR4T g656(.s(BB_361_30110), .d(AA_392), .b(vdd), .g(inst[17]));
NEMR4T g657(.s(BB_361_30110), .d(AA_403), .b(gnd), .g(inst[17]));
NEMR4T g658(.s(BB_361_3011), .d(AA_421), .b(gnd), .g(inst[13]));
NEMR4T g659(.s(BB_361_3011), .d(AA_452), .b(gnd), .g(irq));
NEMR4T g660(.s(next_interrupt_enabled), .d(BB_361_31), .b(gnd), .g(interrupt_enabled));
NEMR4T g661(.s(BB_361_31), .d(BB_361_310), .b(vdd), .g(inst[0]));
NEMR4T g662(.s(BB_361_310), .d(BB_361_3101), .b(gnd), .g(inst[16]));
NEMR4T g663(.s(BB_361_3101), .d(BB_361_31010), .b(vdd), .g(inst[13]));
NEMR4T g664(.s(BB_361_31010), .d(AA_434), .b(vdd), .g(irq));
NEMR4T g665(.s(BB_361_31010), .d(AA_401), .b(gnd), .g(irq));
NEMR4T g666(.s(BB_361_31010), .d(AA_422), .b(vdd), .g(inst[17]));
NEMR4T g667(.s(BB_361_31010), .d(AA_409), .b(gnd), .g(inst[17]));
NEMR4T g668(.s(BB_361_3101), .d(BB_361_31011), .b(gnd), .g(inst[13]));
NEMR4T g669(.s(BB_361_31011), .d(AA_404), .b(gnd), .g(irq));
NEMR4T g670(.s(BB_361_3101), .d(AA_408), .b(gnd), .g(irq));
NEMR4T g671(.s(BB_361_31), .d(BB_361_311), .b(gnd), .g(inst[0]));
NEMR4T g672(.s(BB_361_311), .d(BB_361_3111), .b(gnd), .g(inst[16]));
NEMR4T g673(.s(BB_361_3111), .d(BB_361_31110), .b(vdd), .g(inst[13]));
NEMR4T g674(.s(BB_361_31110), .d(AA_422), .b(vdd), .g(irq));
NEMR4T g675(.s(BB_361_31110), .d(AA_392), .b(gnd), .g(irq));
NEMR4T g676(.s(BB_361_31), .d(BB_361_3120), .b(vdd), .g(inst[16]));
NEMR4T g677(.s(BB_361_3120), .d(AA_435), .b(vdd), .g(irq));
NEMR4T g678(.s(BB_361_3120), .d(AA_392), .b(gnd), .g(irq));
NEMR4T g679(.s(BB_361_31), .d(BB_361_3121), .b(gnd), .g(inst[16]));
NEMR4T g680(.s(BB_361_3121), .d(BB_361_31211), .b(gnd), .g(inst[13]));
NEMR4T g681(.s(BB_361_31211), .d(BB_361_312110), .b(vdd), .g(irq));
NEMR4T g682(.s(BB_361_312110), .d(AA_372), .b(gnd), .g(inst[17]));
NEMR4T g683(.s(AA_372), .d(AA_394), .b(vdd), .g(ireset));
NEMR4T g684(.s(BB_361_312110), .d(AA_392), .b(gnd), .g(ireset));
NEMR4T g685(.s(BB_361_31211), .d(AA_452), .b(gnd), .g(irq));
NEMR4T g686(.s(BB_361_3121), .d(BB_361_312120), .b(vdd), .g(irq));
NEMR4T g687(.s(BB_361_312120), .d(AA_424), .b(vdd), .g(inst[17]));
NEMR4T g688(.s(BB_361_312120), .d(BB_361_3121201), .b(gnd), .g(inst[17]));
NEMR4T g689(.s(BB_361_3121201), .d(AA_391), .b(vdd), .g(ireset));
NEMR4T g690(.s(next_interrupt_enabled), .d(BB_361_321), .b(gnd), .g(inst[0]));
NEMR4T g691(.s(BB_361_321), .d(BB_361_3211), .b(gnd), .g(inst[16]));
NEMR4T g692(.s(BB_361_3211), .d(BB_361_32110), .b(vdd), .g(inst[13]));
NEMR4T g693(.s(BB_361_32110), .d(BB_361_321100), .b(vdd), .g(irq));
NEMR4T g694(.s(BB_361_321100), .d(AA_372), .b(gnd), .g(inst[17]));
NEMR4T g695(.s(BB_361_3211), .d(BB_361_32111), .b(gnd), .g(inst[13]));
NEMR4T g696(.s(BB_361_32111), .d(AA_407), .b(gnd), .g(irq));
NEMR4T g697(.s(werf), .d(BB_373_30), .b(vdd), .g(inst[14]));
NEMR4T g698(.s(BB_373_30), .d(BB_373_300), .b(vdd), .g(inst[16]));
NEMR4T g699(.s(BB_373_300), .d(BB_373_3000), .b(vdd), .g(inst[13]));
NEMR4T g700(.s(BB_373_3000), .d(BB_373_30000), .b(vdd), .g(irq));
NEMR4T g701(.s(BB_373_30000), .d(AA_391), .b(vdd), .g(ireset));
NEMR4T g702(.s(BB_373_30000), .d(AA_395), .b(gnd), .g(ireset));
NEMR4T g703(.s(BB_373_30000), .d(gnd), .b(gnd), .g(inst[15]));
NEMR4T g704(.s(BB_373_3000), .d(AA_392), .b(gnd), .g(irq));
NEMR4T g705(.s(BB_373_30), .d(AA_386), .b(gnd), .g(inst[13]));
NEMR4T g706(.s(AA_386), .d(AA_406), .b(vdd), .g(irq));
NEMR4T g707(.s(AA_386), .d(AA_407), .b(gnd), .g(irq));
NEMR4T g708(.s(AA_386), .d(AA_410), .b(gnd), .g(inst[17]));
NEMR4T g709(.s(werf), .d(BB_373_31), .b(gnd), .g(inst[14]));
NEMR4T g710(.s(BB_373_31), .d(BB_373_310), .b(vdd), .g(inst[16]));
NEMR4T g711(.s(BB_373_310), .d(BB_373_31020), .b(vdd), .g(irq));
NEMR4T g712(.s(BB_373_31020), .d(AA_424), .b(vdd), .g(inst[17]));
NEMR4T g713(.s(BB_373_31020), .d(AA_392), .b(gnd), .g(ireset));
NEMR4T g714(.s(BB_373_310), .d(AA_454), .b(gnd), .g(irq));
NEMR4T g715(.s(BB_373_310), .d(AA_401), .b(gnd), .g(inst[17]));
NEMR4T g716(.s(BB_373_31), .d(BB_373_311), .b(gnd), .g(inst[16]));
NEMR4T g717(.s(BB_373_311), .d(AA_386), .b(gnd), .g(inst[13]));
NEMR4T g718(.s(werf), .d(BB_373_321), .b(gnd), .g(inst[16]));
NEMR4T g719(.s(BB_373_321), .d(AA_386), .b(vdd), .g(inst[13]));
NEMR4T g720(.s(wesp), .d(AA_392), .b(vdd), .g(inst[14]));
NEMR4T g721(.s(wesp), .d(BB_387_31), .b(gnd), .g(inst[14]));
NEMR4T g722(.s(BB_387_31), .d(AA_456), .b(vdd), .g(inst[16]));
NEMR4T g723(.s(BB_387_31), .d(AA_460), .b(gnd), .g(inst[16]));
NEMR4T g724(.s(BB_387_31), .d(AA_392), .b(vdd), .g(inst[13]));
NEMR4T g725(.s(BB_387_31), .d(AA_461), .b(gnd), .g(inst[13]));

endmodule
