module Instruction_decode(clk, ireset, irq, inst, c, z, read_strobe,
     write_strobe, interrupt_ack, next_interrupt_enabled,
     interrupt_enabled, zsel, csel, wsel, pcsel, stsel, werf, wesp);
  input clk, ireset, irq, c, z, interrupt_enabled;
  input [17:0] inst;
  output read_strobe, write_strobe, interrupt_ack,
       next_interrupt_enabled, werf, wesp;
  output [2:0] zsel, csel, wsel;
  output [1:0] pcsel, stsel;

  wire AA_111, AA_117, AA_125, AA_129, AA_136, AA_139, AA_147, AA_148, AA_150, AA_153, 
       AA_154, AA_162, AA_164, AA_165, AA_167, AA_168, AA_169, AA_170, AA_171, AA_173, 
       AA_176, AA_178, AA_179, AA_180, AA_181, AA_182, AA_191, AA_207, AA_214, AA_215, 
       AA_217, AA_220, AA_223, AA_224, AA_225, AA_226, AA_227, AA_228, AA_229, AA_230, 
       AA_231, AA_232, AA_241, AA_242, AA_245, AA_253, AA_260, AA_262, AA_263, AA_264, 
       AA_269, AA_27, AA_272, AA_273, AA_274, AA_275, AA_279, AA_280, AA_281, AA_282, 
       AA_283, AA_284, AA_285, AA_292, AA_294, AA_298, AA_302, AA_308, AA_311, AA_313, 
       AA_325, AA_326, AA_328, AA_334, AA_335, AA_336, AA_340, AA_341, AA_342, AA_372, 
       AA_386, AA_391, AA_392, AA_393, AA_394, AA_395, AA_396, AA_397, AA_398, AA_399, 
       AA_400, AA_401, AA_402, AA_403, AA_404, AA_405, AA_406, AA_407, AA_408, AA_409, 
       AA_410, AA_411, AA_416, AA_419, AA_420, AA_421, AA_422, AA_423, AA_424, AA_425, 
       AA_426, AA_427, AA_428, AA_429, AA_430, AA_431, AA_432, AA_433, AA_434, AA_435, 
       AA_436, AA_441, AA_442, AA_443, AA_444, AA_445, AA_446, AA_447, AA_448, AA_449, 
       AA_450, AA_451, AA_452, AA_453, AA_454, AA_455, AA_456, AA_458, AA_459, AA_460, 
       AA_461, AA_462, AA_463, AA_464, AA_53, AA_79, AA_83, AA_93, BB_0_30, BB_0_3021, 
       BB_0_30211, BB_0_31, BB_0_311, BB_0_3110, BB_0_31100, BB_0_3121, BB_0_320, BB_0_321, BB_0_3211, BB_100_30, 
       BB_100_30222221, BB_100_31, BB_100_310, BB_100_3101, BB_100_31011, BB_100_310221, BB_100_311, BB_100_3110, BB_100_31101, BB_100_311011, 
       BB_100_3111, BB_100_31110, BB_100_31111, BB_100_311111, BB_100_31120, BB_100_31121, BB_100_311211, BB_100_3121, BB_100_31211, BB_100_312110, 
       BB_100_3222220, BB_100_32222201, BB_100_3222221, BB_100_32222211, BB_13_30, BB_13_300, BB_13_3000, BB_13_301, BB_13_3011, BB_13_3021, 
       BB_13_31, BB_13_310, BB_13_320, BB_183_31, BB_183_310, BB_183_3101, BB_183_31011, BB_183_310221, BB_183_311, BB_183_3110, 
       BB_183_31101, BB_183_311011, BB_183_3110111, BB_183_3111, BB_183_31110, BB_183_31111, BB_183_311111, BB_183_3111111, BB_183_31111110, BB_183_311111100, 
       BB_183_31120, BB_183_311201, BB_183_31121, BB_183_311211, BB_183_3112111, BB_183_3121, BB_183_31211, BB_183_312111, BB_183_3121111, BB_233_31, 
       BB_233_310, BB_233_3101, BB_233_31011, BB_233_310221, BB_233_311, BB_233_3110, BB_233_31101, BB_233_311011, BB_233_3111, BB_233_31110, 
       BB_233_31111, BB_233_311111, BB_233_31120, BB_233_31121, BB_233_311211, BB_233_3121, BB_233_31211, BB_286_30, BB_286_30222221, BB_286_31, 
       BB_286_310, BB_286_3101, BB_286_31011, BB_286_310221, BB_286_311, BB_286_3110, BB_286_31101, BB_286_311011, BB_286_3111, BB_286_31110, 
       BB_286_31111, BB_286_311111, BB_286_31120, BB_286_31121, BB_286_311211, BB_286_3121, BB_286_31211, BB_286_312110, BB_286_3222220, BB_286_32222201, 
       BB_286_3222221, BB_286_32222211, BB_28_30, BB_28_301, BB_28_3010, BB_28_31, BB_28_311, BB_28_3111, BB_28_321, BB_28_3211, 
       BB_28_32111, BB_343_31, BB_343_310, BB_343_3100, BB_343_311, BB_343_3121, BB_343_31211, BB_350_30, BB_350_301, BB_350_3010, 
       BB_350_31, BB_350_311, BB_350_321, BB_360_31, BB_361_30, BB_361_301, BB_361_3011, BB_361_30110, BB_361_301100, BB_361_31, 
       BB_361_310, BB_361_3101, BB_361_31010, BB_361_31011, BB_361_311, BB_361_3111, BB_361_31110, BB_361_3120, BB_361_3121, BB_361_31211, 
       BB_361_312110, BB_361_312120, BB_361_3121201, BB_361_321, BB_361_3211, BB_361_32110, BB_361_321100, BB_361_32111, BB_373_30, BB_373_300, 
       BB_373_3000, BB_373_30000, BB_373_31, BB_373_310, BB_373_31020, BB_373_311, BB_373_321, BB_387_31, BB_40_30, BB_40_300, 
       BB_40_31, BB_40_310, BB_40_311, BB_40_3111, BB_40_3121, BB_40_320, BB_40_3201, BB_40_32010, BB_40_32021, BB_40_321, 
       BB_40_3211, BB_40_321220, BB_40_3221, BB_61_30, BB_61_300, BB_61_3000, BB_61_30000, BB_61_31, BB_61_310, BB_61_3101, 
       BB_61_311, BB_61_3110, BB_61_3120, BB_61_320, BB_61_3201, BB_61_32010, BB_61_321, BB_61_3210, BB_61_3211, BB_61_32110, 
       BB_61_321100, BB_61_3220, BB_61_3221, BB_84_30, BB_84_300, BB_84_3000, BB_84_301, BB_84_3010, BB_84_3011, BB_84_31, 
       BB_84_310, BB_84_3101, BB_84_311, BB_84_3111, BB_84_31121, BB_84_320, BB_84_321, BB_84_3210, BB_84_3211, BB_97_30, 
       BB_97_31, BB_97_311, BB_99_31, csel[0], csel[1], csel[2], interrupt_ack, next_interrupt_enabled, pcsel[0], pcsel[1], 
       read_strobe, stsel[0], stsel[1], werf, wesp, write_strobe, wsel[0], wsel[1], zsel[0], zsel[1], zsel[2];

NEMR6T g1(.s1(zsel[0]), .d1(BB_0_30), .s2(zsel[1]), .d2(BB_13_30), .b(vdd), .g(inst[14]));
NEMR6T g2(.s1(BB_0_30), .d1(AA_463), .s2(BB_0_31), .d2(AA_446), .b(vdd), .g(inst[16]));
NEMR6T g3(.s1(AA_463), .d1(AA_458), .s2(BB_0_30), .d2(AA_444), .b(vdd), .g(inst[13]));
NEMR6T g4(.s1(AA_458), .d1(AA_441), .s2(AA_443), .d2(AA_396), .b(vdd), .g(irq));
NEMR6T g5(.s1(AA_441), .d1(AA_391), .s2(AA_444), .d2(AA_398), .b(gnd), .g(inst[17]));
NEMR6T g6(.s1(AA_391), .d1(vdd), .s2(AA_395), .d2(gnd), .b(vdd), .g(inst[15]));
NEMR6T g7(.s1(AA_458), .d1(AA_442), .s2(AA_396), .d2(AA_394), .b(vdd), .g(inst[17]));
NEMR6T g8(.s1(AA_442), .d1(AA_392), .s2(AA_396), .d2(AA_395), .b(vdd), .g(ireset));
NEMR6T g9(.s1(AA_392), .d1(gnd), .s2(AA_393), .d2(vdd), .b(gnd), .g(vdd));
NEMR6T g10(.s1(AA_442), .d1(AA_393), .s2(AA_396), .d2(AA_391), .b(gnd), .g(ireset));
NEMR6T g11(.s1(BB_0_30), .d1(AA_443), .s2(BB_0_31), .d2(BB_0_311), .b(gnd), .g(inst[16]));
NEMR6T g12(.s1(AA_394), .d1(vdd), .s2(AA_397), .d2(gnd), .b(gnd), .g(inst[15]));
NEMR6T g13(.s1(AA_398), .d1(AA_397), .s2(AA_399), .d2(AA_395), .b(vdd), .g(ireset));
NEMR6T g14(.s1(AA_398), .d1(AA_394), .s2(AA_399), .d2(AA_391), .b(gnd), .g(ireset));
NEMR6T g15(.s1(BB_0_30), .d1(BB_0_3021), .s2(BB_0_311), .d2(AA_443), .b(gnd), .g(inst[13]));
NEMR6T g16(.s1(BB_0_3021), .d1(BB_0_30211), .s2(BB_0_30), .d2(AA_445), .b(gnd), .g(irq));
NEMR6T g17(.s1(BB_0_30211), .d1(AA_442), .s2(BB_0_31100), .d2(AA_393), .b(vdd), .g(inst[17]));
NEMR6T g18(.s1(BB_0_30211), .d1(AA_398), .s2(AA_445), .d2(AA_399), .b(gnd), .g(inst[17]));
NEMR6T g19(.s1(zsel[0]), .d1(BB_0_31), .s2(zsel[1]), .d2(BB_13_31), .b(gnd), .g(inst[14]));
NEMR6T g20(.s1(AA_446), .d1(AA_442), .s2(BB_0_311), .d2(BB_0_3110), .b(vdd), .g(inst[13]));
NEMR6T g21(.s1(BB_0_3110), .d1(BB_0_31100), .s2(AA_447), .d2(AA_442), .b(vdd), .g(irq));
NEMR6T g22(.s1(BB_0_3110), .d1(AA_442), .s2(AA_449), .d2(AA_400), .b(gnd), .g(inst[17]));
NEMR6T g23(.s1(BB_0_31), .d1(BB_0_3121), .s2(BB_0_320), .d2(AA_447), .b(gnd), .g(inst[13]));
NEMR6T g24(.s1(BB_0_3121), .d1(AA_442), .s2(AA_459), .d2(AA_448), .b(gnd), .g(irq));
NEMR6T g25(.s1(zsel[0]), .d1(BB_0_320), .s2(BB_13_30), .d2(BB_13_300), .b(vdd), .g(inst[16]));
NEMR6T g26(.s1(zsel[0]), .d1(BB_0_321), .s2(BB_13_30), .d2(BB_13_301), .b(gnd), .g(inst[16]));
NEMR6T g27(.s1(BB_0_321), .d1(AA_459), .s2(BB_13_300), .d2(BB_13_3000), .b(vdd), .g(inst[13]));
NEMR6T g28(.s1(AA_448), .d1(AA_442), .s2(BB_13_3000), .d2(AA_392), .b(vdd), .g(inst[17]));
NEMR6T g29(.s1(BB_0_321), .d1(BB_0_3211), .s2(BB_13_301), .d2(BB_13_3011), .b(gnd), .g(inst[13]));
NEMR6T g30(.s1(BB_0_3211), .d1(AA_444), .s2(BB_13_3000), .d2(AA_449), .b(vdd), .g(irq));
NEMR6T g31(.s1(AA_400), .d1(AA_391), .s2(AA_401), .d2(AA_392), .b(vdd), .g(ireset));
NEMR6T g32(.s1(AA_400), .d1(gnd), .s2(BB_99_31), .d2(gnd), .b(gnd), .g(inst[15]));
NEMR6T g33(.s1(BB_13_300), .d1(AA_450), .s2(BB_13_3021), .d2(AA_404), .b(gnd), .g(irq));
NEMR6T g34(.s1(AA_450), .d1(AA_401), .s2(BB_13_3011), .d2(AA_403), .b(gnd), .g(inst[17]));
NEMR6T g35(.s1(BB_13_3011), .d1(AA_402), .s2(BB_13_3021), .d2(AA_450), .b(vdd), .g(irq));
NEMR6T g36(.s1(AA_402), .d1(AA_400), .s2(AA_404), .d2(AA_392), .b(vdd), .g(inst[17]));
NEMR6T g37(.s1(AA_402), .d1(AA_395), .s2(AA_403), .d2(AA_397), .b(gnd), .g(ireset));
NEMR6T g38(.s1(BB_13_30), .d1(BB_13_3021), .s2(AA_460), .d2(AA_451), .b(gnd), .g(inst[13]));
NEMR6T g39(.s1(BB_13_31), .d1(BB_13_310), .s2(zsel[1]), .d2(BB_13_320), .b(vdd), .g(inst[16]));
NEMR6T g40(.s1(BB_13_310), .d1(AA_27), .s2(AA_464), .d2(AA_392), .b(vdd), .g(inst[13]));
NEMR6T g41(.s1(AA_27), .d1(AA_406), .s2(AA_451), .d2(AA_392), .b(vdd), .g(irq));
NEMR6T g42(.s1(AA_406), .d1(AA_405), .s2(AA_407), .d2(AA_392), .b(vdd), .g(inst[17]));
NEMR6T g43(.s1(AA_405), .d1(AA_394), .s2(AA_410), .d2(AA_392), .b(vdd), .g(ireset));
NEMR6T g44(.s1(AA_405), .d1(gnd), .s2(BB_99_31), .d2(vdd), .b(vdd), .g(inst[15]));
NEMR6T g45(.s1(AA_406), .d1(AA_397), .s2(AA_409), .d2(AA_395), .b(gnd), .g(ireset));
NEMR6T g46(.s1(BB_13_310), .d1(AA_404), .s2(AA_451), .d2(AA_407), .b(gnd), .g(irq));
NEMR6T g47(.s1(BB_13_310), .d1(AA_401), .s2(AA_407), .d2(AA_403), .b(gnd), .g(inst[17]));
NEMR6T g48(.s1(BB_13_31), .d1(AA_460), .s2(zsel[1]), .d2(AA_464), .b(gnd), .g(inst[16]));
NEMR6T g49(.s1(BB_13_320), .d1(AA_27), .s2(AA_464), .d2(AA_461), .b(gnd), .g(inst[13]));
NEMR6T g50(.s1(BB_13_320), .d1(AA_408), .s2(AA_461), .d2(AA_452), .b(gnd), .g(irq));
NEMR6T g51(.s1(AA_408), .d1(AA_403), .s2(BB_13_320), .d2(AA_409), .b(gnd), .g(inst[17]));
NEMR6T g52(.s1(AA_452), .d1(AA_410), .s2(AA_411), .d2(AA_394), .b(gnd), .g(inst[17]));
NEMR6T g53(.s1(AA_410), .d1(AA_395), .s2(BB_61_321100), .d2(AA_394), .b(gnd), .g(ireset));
NEMR6T g54(.s1(zsel[2]), .d1(BB_28_30), .s2(BB_40_30), .d2(BB_40_300), .b(vdd), .g(inst[14]));
NEMR6T g55(.s1(BB_28_30), .d1(BB_28_301), .s2(BB_28_31), .d2(BB_28_311), .b(gnd), .g(inst[16]));
NEMR6T g56(.s1(BB_28_301), .d1(BB_28_3010), .s2(BB_28_311), .d2(AA_442), .b(vdd), .g(inst[13]));
NEMR6T g57(.s1(BB_28_3010), .d1(AA_411), .s2(BB_28_3211), .d2(AA_442), .b(vdd), .g(irq));
NEMR6T g58(.s1(BB_28_3010), .d1(AA_442), .s2(BB_28_32111), .d2(AA_442), .b(vdd), .g(inst[17]));
NEMR6T g59(.s1(BB_28_3010), .d1(AA_399), .s2(BB_28_32111), .d2(AA_399), .b(gnd), .g(inst[17]));
NEMR6T g60(.s1(BB_28_301), .d1(AA_444), .s2(BB_28_3111), .d2(AA_444), .b(gnd), .g(irq));
NEMR6T g61(.s1(zsel[2]), .d1(BB_28_31), .s2(BB_40_30), .d2(AA_416), .b(gnd), .g(inst[14]));
NEMR6T g62(.s1(BB_28_311), .d1(BB_28_3111), .s2(BB_28_321), .d2(BB_28_3211), .b(gnd), .g(inst[13]));
NEMR6T g63(.s1(zsel[2]), .d1(AA_442), .s2(BB_40_300), .d2(AA_446), .b(vdd), .g(inst[16]));
NEMR6T g64(.s1(zsel[2]), .d1(BB_28_321), .s2(BB_40_311), .d2(BB_40_3111), .b(gnd), .g(inst[16]));
NEMR6T g65(.s1(BB_28_3211), .d1(BB_28_32111), .s2(AA_416), .d2(AA_445), .b(gnd), .g(irq));
NEMR6T g66(.s1(csel[0]), .d1(BB_40_30), .s2(csel[1]), .d2(BB_61_30), .b(vdd), .g(inst[3]));
NEMR6T g67(.s1(BB_40_300), .d1(AA_416), .s2(BB_40_3121), .d2(AA_416), .b(gnd), .g(inst[13]));
NEMR6T g68(.s1(AA_416), .d1(AA_398), .s2(BB_84_3000), .d2(AA_409), .b(gnd), .g(inst[17]));
NEMR6T g69(.s1(csel[0]), .d1(BB_40_31), .s2(csel[1]), .d2(BB_61_31), .b(gnd), .g(inst[3]));
NEMR6T g70(.s1(BB_40_31), .d1(BB_40_310), .s2(csel[0]), .d2(BB_40_320), .b(vdd), .g(inst[14]));
NEMR6T g71(.s1(BB_40_310), .d1(AA_463), .s2(BB_40_31), .d2(AA_416), .b(vdd), .g(inst[16]));
NEMR6T g72(.s1(BB_40_31), .d1(BB_40_311), .s2(csel[0]), .d2(BB_40_321), .b(gnd), .g(inst[14]));
NEMR6T g73(.s1(BB_40_3111), .d1(AA_416), .s2(BB_40_3201), .d2(BB_40_32010), .b(vdd), .g(inst[13]));
NEMR6T g74(.s1(BB_40_31), .d1(BB_40_3121), .s2(BB_40_320), .d2(BB_40_3201), .b(gnd), .g(inst[16]));
NEMR6T g75(.s1(BB_40_32010), .d1(AA_394), .s2(BB_40_32021), .d2(AA_396), .b(vdd), .g(irq));
NEMR6T g76(.s1(BB_40_32010), .d1(AA_442), .s2(BB_40_32021), .d2(AA_448), .b(gnd), .g(irq));
NEMR6T g77(.s1(BB_40_320), .d1(BB_40_32021), .s2(BB_40_3211), .d2(AA_53), .b(gnd), .g(inst[13]));
NEMR6T g78(.s1(BB_40_321), .d1(AA_53), .s2(BB_61_300), .d2(BB_61_3000), .b(vdd), .g(inst[16]));
NEMR6T g79(.s1(AA_53), .d1(AA_399), .s2(BB_40_321), .d2(BB_40_321220), .b(vdd), .g(irq));
NEMR6T g80(.s1(BB_40_321), .d1(BB_40_3211), .s2(csel[0]), .d2(BB_40_3221), .b(gnd), .g(inst[16]));
NEMR6T g81(.s1(BB_40_321220), .d1(AA_394), .s2(BB_61_321100), .d2(AA_391), .b(vdd), .g(inst[17]));
NEMR6T g82(.s1(BB_40_321), .d1(AA_448), .s2(AA_79), .d2(AA_445), .b(gnd), .g(irq));
NEMR6T g83(.s1(BB_40_3221), .d1(AA_53), .s2(BB_61_3000), .d2(BB_61_30000), .b(vdd), .g(inst[13]));
NEMR6T g84(.s1(BB_61_30), .d1(BB_61_300), .s2(BB_61_31), .d2(BB_61_310), .b(vdd), .g(inst[14]));
NEMR6T g85(.s1(BB_61_30000), .d1(AA_441), .s2(BB_61_32010), .d2(AA_411), .b(vdd), .g(irq));
NEMR6T g86(.s1(BB_61_300), .d1(AA_448), .s2(BB_61_3101), .d2(AA_448), .b(vdd), .g(inst[13]));
NEMR6T g87(.s1(BB_61_30), .d1(AA_416), .s2(BB_61_310), .d2(AA_446), .b(vdd), .g(inst[16]));
NEMR6T g88(.s1(BB_61_30), .d1(AA_83), .s2(BB_61_310), .d2(BB_61_3101), .b(gnd), .g(inst[16]));
NEMR6T g89(.s1(AA_83), .d1(AA_79), .s2(BB_61_310), .d2(AA_79), .b(gnd), .g(inst[13]));
NEMR6T g90(.s1(BB_61_31), .d1(BB_61_311), .s2(csel[1]), .d2(BB_61_321), .b(gnd), .g(inst[14]));
NEMR6T g91(.s1(BB_61_311), .d1(BB_61_3110), .s2(BB_61_31), .d2(BB_61_3120), .b(vdd), .g(inst[16]));
NEMR6T g92(.s1(BB_61_3110), .d1(AA_444), .s2(BB_61_3201), .d2(BB_61_32010), .b(vdd), .g(inst[13]));
NEMR6T g93(.s1(BB_61_3110), .d1(AA_445), .s2(BB_61_321), .d2(AA_448), .b(gnd), .g(irq));
NEMR6T g94(.s1(BB_61_311), .d1(AA_83), .s2(BB_61_320), .d2(BB_61_3201), .b(gnd), .g(inst[16]));
NEMR6T g95(.s1(BB_61_3120), .d1(AA_444), .s2(BB_61_320), .d2(AA_459), .b(gnd), .g(inst[13]));
NEMR6T g96(.s1(csel[1]), .d1(BB_61_320), .s2(csel[2]), .d2(BB_84_30), .b(vdd), .g(inst[14]));
NEMR6T g97(.s1(BB_61_321), .d1(BB_61_3210), .s2(csel[1]), .d2(BB_61_3220), .b(vdd), .g(inst[16]));
NEMR6T g98(.s1(BB_61_3210), .d1(AA_443), .s2(BB_61_3211), .d2(BB_61_32110), .b(vdd), .g(inst[13]));
NEMR6T g99(.s1(BB_61_321), .d1(BB_61_3211), .s2(csel[1]), .d2(BB_61_3221), .b(gnd), .g(inst[16]));
NEMR6T g100(.s1(BB_61_32110), .d1(BB_61_321100), .s2(BB_84_3000), .d2(AA_449), .b(vdd), .g(irq));
NEMR6T g101(.s1(BB_61_321100), .d1(AA_397), .s2(AA_423), .d2(AA_392), .b(vdd), .g(ireset));
NEMR6T g102(.s1(BB_61_3220), .d1(AA_443), .s2(BB_61_3221), .d2(AA_447), .b(gnd), .g(inst[13]));
NEMR6T g103(.s1(BB_61_3221), .d1(AA_445), .s2(BB_84_300), .d2(BB_84_3000), .b(vdd), .g(inst[13]));
NEMR6T g104(.s1(BB_61_3221), .d1(AA_444), .s2(BB_84_300), .d2(AA_408), .b(gnd), .g(irq));
NEMR6T g105(.s1(BB_84_30), .d1(BB_84_300), .s2(BB_84_31), .d2(BB_84_310), .b(vdd), .g(inst[16]));
NEMR6T g106(.s1(BB_84_30), .d1(BB_84_301), .s2(BB_84_31), .d2(BB_84_311), .b(gnd), .g(inst[16]));
NEMR6T g107(.s1(BB_84_301), .d1(BB_84_3010), .s2(BB_84_30), .d2(AA_404), .b(vdd), .g(inst[13]));
NEMR6T g108(.s1(BB_84_3010), .d1(AA_419), .s2(BB_84_3011), .d2(AA_402), .b(vdd), .g(irq));
NEMR6T g109(.s1(AA_419), .d1(AA_405), .s2(BB_84_301), .d2(AA_403), .b(gnd), .g(inst[17]));
NEMR6T g110(.s1(BB_84_301), .d1(BB_84_3011), .s2(BB_84_30), .d2(AA_453), .b(gnd), .g(inst[13]));
NEMR6T g111(.s1(AA_453), .d1(AA_420), .s2(BB_84_30), .d2(AA_450), .b(gnd), .g(irq));
NEMR6T g112(.s1(AA_420), .d1(AA_392), .s2(AA_454), .d2(AA_392), .b(vdd), .g(inst[17]));
NEMR6T g113(.s1(AA_420), .d1(AA_409), .s2(AA_454), .d2(AA_422), .b(gnd), .g(inst[17]));
NEMR6T g114(.s1(csel[2]), .d1(BB_84_31), .s2(wsel[0]), .d2(BB_97_31), .b(gnd), .g(inst[14]));
NEMR6T g115(.s1(BB_84_310), .d1(AA_392), .s2(BB_84_311), .d2(AA_421), .b(vdd), .g(inst[13]));
NEMR6T g116(.s1(BB_84_310), .d1(BB_84_3101), .s2(BB_84_311), .d2(BB_84_3111), .b(gnd), .g(inst[13]));
NEMR6T g117(.s1(BB_84_3101), .d1(AA_392), .s2(BB_84_3111), .d2(AA_93), .b(gnd), .g(irq));
NEMR6T g118(.s1(AA_421), .d1(AA_392), .s2(BB_84_3111), .d2(AA_454), .b(vdd), .g(irq));
NEMR6T g119(.s1(AA_422), .d1(AA_392), .s2(AA_423), .d2(AA_397), .b(gnd), .g(ireset));
NEMR6T g120(.s1(AA_93), .d1(AA_409), .s2(BB_84_31121), .d2(AA_423), .b(gnd), .g(inst[17]));
NEMR6T g121(.s1(BB_84_311), .d1(BB_84_31121), .s2(BB_84_3210), .d2(AA_93), .b(gnd), .g(irq));
NEMR6T g122(.s1(BB_84_31121), .d1(AA_392), .s2(BB_97_30), .d2(AA_392), .b(vdd), .g(inst[17]));
NEMR6T g123(.s1(csel[2]), .d1(BB_84_320), .s2(AA_179), .d2(AA_178), .b(vdd), .g(inst[16]));
NEMR6T g124(.s1(BB_84_320), .d1(AA_421), .s2(BB_84_321), .d2(BB_84_3211), .b(gnd), .g(inst[13]));
NEMR6T g125(.s1(csel[2]), .d1(BB_84_321), .s2(AA_182), .d2(AA_180), .b(gnd), .g(inst[16]));
NEMR6T g126(.s1(BB_84_321), .d1(BB_84_3210), .s2(BB_97_31), .d2(AA_391), .b(vdd), .g(inst[13]));
NEMR6T g127(.s1(BB_84_3211), .d1(AA_450), .s2(AA_167), .d2(AA_411), .b(vdd), .g(irq));
NEMR6T g128(.s1(wsel[0]), .d1(BB_97_30), .s2(wsel[1]), .d2(AA_392), .b(vdd), .g(inst[14]));
NEMR6T g129(.s1(BB_97_30), .d1(AA_393), .s2(BB_97_311), .d2(AA_391), .b(gnd), .g(inst[17]));
NEMR6T g130(.s1(BB_97_31), .d1(BB_97_311), .s2(AA_178), .d2(AA_167), .b(gnd), .g(inst[13]));
NEMR6T g131(.s1(BB_97_311), .d1(AA_395), .s2(BB_97_31), .d2(AA_397), .b(vdd), .g(inst[17]));
NEMR6T g132(.s1(BB_97_31), .d1(AA_394), .s2(AA_167), .d2(AA_426), .b(gnd), .g(inst[17]));
NEMR6T g133(.s1(wsel[1]), .d1(BB_99_31), .s2(BB_100_30), .d2(AA_182), .b(gnd), .g(inst[14]));
NEMR6T g134(.s1(pcsel[1]), .d1(BB_100_30), .s2(pcsel[0]), .d2(AA_231), .b(vdd), .g(inst[12]));
NEMR6T g135(.s1(BB_100_30), .d1(AA_179), .s2(AA_173), .d2(AA_154), .b(vdd), .g(inst[14]));
NEMR6T g136(.s1(AA_167), .d1(AA_424), .s2(AA_169), .d2(AA_147), .b(gnd), .g(irq));
NEMR6T g137(.s1(AA_424), .d1(AA_393), .s2(AA_427), .d2(AA_395), .b(vdd), .g(ireset));
NEMR6T g138(.s1(AA_167), .d1(AA_425), .s2(AA_168), .d2(AA_401), .b(vdd), .g(inst[17]));
NEMR6T g139(.s1(AA_425), .d1(AA_393), .s2(AA_426), .d2(AA_391), .b(gnd), .g(ireset));
NEMR6T g140(.s1(AA_179), .d1(AA_169), .s2(AA_148), .d2(AA_429), .b(gnd), .g(inst[13]));
NEMR6T g141(.s1(AA_169), .d1(AA_168), .s2(AA_429), .d2(AA_442), .b(vdd), .g(irq));
NEMR6T g142(.s1(AA_168), .d1(AA_427), .s2(AA_147), .d2(AA_428), .b(gnd), .g(inst[17]));
NEMR6T g143(.s1(AA_428), .d1(AA_394), .s2(AA_111), .d2(AA_391), .b(gnd), .g(ireset));
NEMR6T g144(.s1(AA_182), .d1(AA_148), .s2(BB_100_30), .d2(AA_431), .b(vdd), .g(inst[16]));
NEMR6T g145(.s1(AA_429), .d1(AA_393), .s2(AA_171), .d2(AA_150), .b(gnd), .g(irq));
NEMR6T g146(.s1(AA_180), .d1(AA_171), .s2(AA_431), .d2(AA_429), .b(vdd), .g(inst[13]));
NEMR6T g147(.s1(AA_171), .d1(AA_170), .s2(AA_153), .d2(AA_117), .b(vdd), .g(irq));
NEMR6T g148(.s1(AA_170), .d1(AA_430), .s2(AA_150), .d2(AA_111), .b(gnd), .g(inst[17]));
NEMR6T g149(.s1(AA_430), .d1(AA_397), .s2(AA_111), .d2(AA_393), .b(vdd), .g(ireset));
NEMR6T g150(.s1(AA_150), .d1(AA_393), .s2(AA_224), .d2(AA_425), .b(vdd), .g(inst[17]));
NEMR6T g151(.s1(BB_100_30), .d1(BB_100_30222221), .s2(AA_154), .d2(AA_169), .b(gnd), .g(inst[16]));
NEMR6T g152(.s1(BB_100_30222221), .d1(AA_169), .s2(AA_455), .d2(AA_432), .b(vdd), .g(inst[13]));
NEMR6T g153(.s1(BB_100_30222221), .d1(AA_153), .s2(AA_164), .d2(AA_153), .b(gnd), .g(inst[13]));
NEMR6T g154(.s1(AA_117), .d1(AA_430), .s2(AA_224), .d2(AA_428), .b(gnd), .g(inst[17]));
NEMR6T g155(.s1(AA_117), .d1(AA_393), .s2(AA_214), .d2(AA_393), .b(gnd), .g(ireset));
NEMR6T g156(.s1(AA_153), .d1(AA_150), .s2(AA_432), .d2(AA_393), .b(gnd), .g(irq));
NEMR6T g157(.s1(pcsel[1]), .d1(BB_100_31), .s2(pcsel[0]), .d2(BB_183_31), .b(gnd), .g(inst[12]));
NEMR6T g158(.s1(BB_100_31), .d1(BB_100_310), .s2(BB_183_31), .d2(BB_183_310), .b(vdd), .g(z));
NEMR6T g159(.s1(BB_100_310), .d1(AA_181), .s2(BB_100_311), .d2(BB_100_3110), .b(vdd), .g(c));
NEMR6T g160(.s1(AA_181), .d1(AA_173), .s2(BB_100_31101), .d2(AA_173), .b(vdd), .g(inst[10]));
NEMR6T g161(.s1(AA_173), .d1(AA_462), .s2(BB_100_310221), .d2(AA_182), .b(gnd), .g(inst[14]));
NEMR6T g162(.s1(AA_462), .d1(AA_455), .s2(AA_176), .d2(AA_125), .b(gnd), .g(inst[16]));
NEMR6T g163(.s1(AA_432), .d1(AA_401), .s2(AA_433), .d2(AA_425), .b(vdd), .g(irq));
NEMR6T g164(.s1(AA_173), .d1(AA_429), .s2(AA_176), .d2(AA_431), .b(vdd), .g(inst[16]));
NEMR6T g165(.s1(AA_181), .d1(AA_176), .s2(BB_100_31011), .d2(AA_162), .b(gnd), .g(inst[10]));
NEMR6T g166(.s1(AA_176), .d1(AA_179), .s2(AA_162), .d2(AA_129), .b(vdd), .g(inst[14]));
NEMR6T g167(.s1(AA_125), .d1(AA_169), .s2(BB_100_32222201), .d2(AA_167), .b(vdd), .g(inst[13]));
NEMR6T g168(.s1(BB_100_310), .d1(BB_100_3101), .s2(BB_100_311), .d2(BB_100_3111), .b(gnd), .g(c));
NEMR6T g169(.s1(BB_100_3101), .d1(AA_181), .s2(BB_100_3111), .d2(BB_100_31110), .b(vdd), .g(inst[11]));
NEMR6T g170(.s1(BB_100_3101), .d1(BB_100_31011), .s2(BB_100_3110), .d2(BB_100_31101), .b(gnd), .g(inst[11]));
NEMR6T g171(.s1(AA_129), .d1(AA_429), .s2(AA_136), .d2(AA_431), .b(vdd), .g(inst[16]));
NEMR6T g172(.s1(AA_129), .d1(AA_169), .s2(BB_100_310), .d2(AA_164), .b(gnd), .g(inst[16]));
NEMR6T g173(.s1(BB_100_310), .d1(BB_100_310221), .s2(BB_100_31101), .d2(BB_100_311011), .b(gnd), .g(inst[10]));
NEMR6T g174(.s1(BB_100_31), .d1(BB_100_311), .s2(BB_183_31), .d2(BB_183_311), .b(gnd), .g(z));
NEMR6T g175(.s1(BB_100_311011), .d1(AA_179), .s2(BB_100_311111), .d2(AA_148), .b(vdd), .g(inst[14]));
NEMR6T g176(.s1(BB_100_3110), .d1(AA_165), .s2(BB_100_31110), .d2(AA_165), .b(gnd), .g(inst[10]));
NEMR6T g177(.s1(AA_165), .d1(AA_136), .s2(BB_100_311111), .d2(AA_139), .b(gnd), .g(inst[14]));
NEMR6T g178(.s1(AA_136), .d1(AA_125), .s2(BB_100_3110), .d2(AA_164), .b(gnd), .g(inst[16]));
NEMR6T g179(.s1(BB_100_31110), .d1(AA_164), .s2(AA_139), .d2(AA_164), .b(gnd), .g(inst[16]));
NEMR6T g180(.s1(BB_100_3111), .d1(BB_100_31111), .s2(BB_100_311), .d2(BB_100_31121), .b(gnd), .g(inst[11]));
NEMR6T g181(.s1(BB_100_31111), .d1(AA_139), .s2(BB_100_31120), .d2(AA_176), .b(vdd), .g(inst[10]));
NEMR6T g182(.s1(BB_100_31111), .d1(BB_100_311111), .s2(BB_100_31120), .d2(AA_162), .b(gnd), .g(inst[10]));
NEMR6T g183(.s1(BB_100_311), .d1(BB_100_31120), .s2(BB_183_3101), .d2(AA_232), .b(vdd), .g(inst[11]));
NEMR6T g184(.s1(BB_100_31120), .d1(AA_182), .s2(BB_100_311211), .d2(AA_182), .b(gnd), .g(inst[14]));
NEMR6T g185(.s1(BB_100_31121), .d1(BB_100_311211), .s2(BB_100_31211), .d2(AA_165), .b(gnd), .g(inst[10]));
NEMR6T g186(.s1(BB_100_311211), .d1(AA_136), .s2(BB_100_312110), .d2(AA_179), .b(vdd), .g(inst[14]));
NEMR6T g187(.s1(BB_100_31), .d1(BB_100_3121), .s2(BB_183_310), .d2(BB_183_3101), .b(gnd), .g(c));
NEMR6T g188(.s1(BB_100_3121), .d1(BB_100_31211), .s2(BB_183_3101), .d2(BB_183_31011), .b(gnd), .g(inst[11]));
NEMR6T g189(.s1(BB_100_31211), .d1(BB_100_312110), .s2(AA_232), .d2(AA_429), .b(vdd), .g(inst[10]));
NEMR6T g190(.s1(BB_100_312110), .d1(AA_182), .s2(pcsel[1]), .d2(BB_100_3222221), .b(gnd), .g(inst[14]));
NEMR6T g191(.s1(BB_100_312110), .d1(AA_431), .s2(AA_231), .d2(AA_429), .b(vdd), .g(inst[16]));
NEMR6T g192(.s1(BB_100_312110), .d1(AA_125), .s2(BB_100_3222220), .d2(BB_100_32222201), .b(gnd), .g(inst[16]));
NEMR6T g193(.s1(pcsel[1]), .d1(BB_100_3222220), .s2(AA_284), .d2(AA_280), .b(vdd), .g(inst[14]));
NEMR6T g194(.s1(BB_100_3222221), .d1(BB_100_32222211), .s2(AA_231), .d2(AA_227), .b(gnd), .g(inst[16]));
NEMR6T g195(.s1(BB_100_32222211), .d1(AA_433), .s2(AA_227), .d2(AA_224), .b(vdd), .g(inst[13]));
NEMR6T g196(.s1(BB_100_32222211), .d1(AA_169), .s2(AA_227), .d2(AA_225), .b(gnd), .g(inst[13]));
NEMR6T g197(.s1(AA_224), .d1(AA_441), .s2(AA_225), .d2(AA_214), .b(vdd), .g(irq));
NEMR6T g198(.s1(AA_224), .d1(AA_424), .s2(AA_225), .d2(AA_215), .b(gnd), .g(irq));
NEMR6T g199(.s1(AA_214), .d1(AA_427), .s2(AA_215), .d2(AA_191), .b(gnd), .g(inst[17]));
NEMR6T g200(.s1(AA_215), .d1(AA_393), .s2(AA_226), .d2(AA_401), .b(vdd), .g(inst[17]));
NEMR6T g201(.s1(AA_191), .d1(AA_393), .s2(AA_260), .d2(AA_391), .b(vdd), .g(ireset));
NEMR6T g202(.s1(AA_191), .d1(AA_394), .s2(AA_260), .d2(AA_395), .b(gnd), .g(ireset));
NEMR6T g203(.s1(AA_227), .d1(AA_226), .s2(AA_220), .d2(AA_226), .b(vdd), .g(irq));
NEMR6T g204(.s1(AA_226), .d1(AA_430), .s2(AA_217), .d2(AA_426), .b(gnd), .g(inst[17]));
NEMR6T g205(.s1(AA_227), .d1(AA_217), .s2(AA_220), .d2(AA_217), .b(gnd), .g(irq));
NEMR6T g206(.s1(BB_183_310), .d1(AA_232), .s2(BB_183_311), .d2(BB_183_3110), .b(vdd), .g(c));
NEMR6T g207(.s1(AA_232), .d1(AA_228), .s2(BB_183_31011), .d2(AA_462), .b(gnd), .g(inst[10]));
NEMR6T g208(.s1(AA_228), .d1(AA_220), .s2(BB_183_310221), .d2(AA_229), .b(gnd), .g(inst[16]));
NEMR6T g209(.s1(AA_220), .d1(AA_224), .s2(BB_183_3110111), .d2(AA_224), .b(vdd), .g(inst[13]));
NEMR6T g210(.s1(BB_183_310), .d1(BB_183_310221), .s2(BB_183_31101), .d2(BB_183_311011), .b(gnd), .g(inst[10]));
NEMR6T g211(.s1(BB_183_310221), .d1(AA_429), .s2(BB_183_31120), .d2(AA_429), .b(vdd), .g(inst[16]));
NEMR6T g212(.s1(AA_229), .d1(AA_225), .s2(AA_223), .d2(AA_207), .b(gnd), .g(inst[13]));
NEMR6T g213(.s1(BB_183_3110), .d1(BB_183_31101), .s2(BB_183_3111), .d2(BB_183_31111), .b(gnd), .g(inst[11]));
NEMR6T g214(.s1(BB_183_31101), .d1(AA_429), .s2(BB_183_31120), .d2(AA_228), .b(vdd), .g(inst[10]));
NEMR6T g215(.s1(BB_183_311011), .d1(BB_183_3110111), .s2(AA_230), .d2(AA_223), .b(gnd), .g(inst[16]));
NEMR6T g216(.s1(BB_183_3110), .d1(AA_230), .s2(BB_183_31110), .d2(AA_230), .b(gnd), .g(inst[10]));
NEMR6T g217(.s1(AA_207), .d1(AA_226), .s2(BB_183_31111110), .d2(BB_183_311111100), .b(vdd), .g(irq));
NEMR6T g218(.s1(AA_207), .d1(AA_217), .s2(BB_183_31111110), .d2(AA_215), .b(gnd), .g(irq));
NEMR6T g219(.s1(BB_183_311), .d1(BB_183_3111), .s2(BB_183_31), .d2(BB_183_3121), .b(gnd), .g(c));
NEMR6T g220(.s1(BB_183_3111), .d1(BB_183_31110), .s2(BB_183_311), .d2(BB_183_31120), .b(vdd), .g(inst[11]));
NEMR6T g221(.s1(BB_183_31111), .d1(BB_183_311111), .s2(BB_183_31120), .d2(BB_183_311201), .b(gnd), .g(inst[10]));
NEMR6T g222(.s1(BB_183_311111), .d1(BB_183_3111111), .s2(BB_183_311201), .d2(AA_431), .b(gnd), .g(inst[16]));
NEMR6T g223(.s1(BB_183_3111111), .d1(BB_183_31111110), .s2(BB_183_3112111), .d2(AA_207), .b(vdd), .g(inst[13]));
NEMR6T g224(.s1(BB_183_311111100), .d1(AA_427), .s2(AA_434), .d2(AA_397), .b(gnd), .g(inst[17]));
NEMR6T g225(.s1(BB_183_31120), .d1(AA_229), .s2(BB_183_311211), .d2(BB_183_3112111), .b(gnd), .g(inst[16]));
NEMR6T g226(.s1(BB_183_311), .d1(BB_183_31121), .s2(BB_183_3121), .d2(BB_183_31211), .b(gnd), .g(inst[11]));
NEMR6T g227(.s1(BB_183_31121), .d1(BB_183_311211), .s2(BB_183_31211), .d2(BB_183_312111), .b(gnd), .g(inst[10]));
NEMR6T g228(.s1(BB_183_311211), .d1(AA_429), .s2(AA_284), .d2(AA_242), .b(vdd), .g(inst[16]));
NEMR6T g229(.s1(BB_183_3112111), .d1(AA_225), .s2(BB_183_3121111), .d2(AA_207), .b(gnd), .g(inst[13]));
NEMR6T g230(.s1(BB_183_31211), .d1(AA_231), .s2(AA_285), .d2(AA_242), .b(vdd), .g(inst[10]));
NEMR6T g231(.s1(BB_183_312111), .d1(BB_183_3121111), .s2(AA_280), .d2(AA_273), .b(gnd), .g(inst[16]));
NEMR6T g232(.s1(BB_183_3121111), .d1(AA_433), .s2(AA_273), .d2(AA_272), .b(vdd), .g(inst[13]));
NEMR6T g233(.s1(stsel[0]), .d1(AA_284), .s2(stsel[1]), .d2(BB_286_30), .b(vdd), .g(inst[12]));
NEMR6T g234(.s1(AA_272), .d1(AA_434), .s2(AA_273), .d2(AA_404), .b(vdd), .g(irq));
NEMR6T g235(.s1(AA_272), .d1(AA_260), .s2(AA_262), .d2(AA_241), .b(gnd), .g(inst[17]));
NEMR6T g236(.s1(AA_273), .d1(AA_262), .s2(AA_242), .d2(AA_435), .b(gnd), .g(irq));
NEMR6T g237(.s1(AA_262), .d1(AA_435), .s2(AA_436), .d2(AA_392), .b(vdd), .g(inst[17]));
NEMR6T g238(.s1(AA_435), .d1(AA_393), .s2(AA_241), .d2(AA_394), .b(vdd), .g(ireset));
NEMR6T g239(.s1(AA_435), .d1(AA_392), .s2(AA_241), .d2(AA_397), .b(gnd), .g(ireset));
NEMR6T g240(.s1(AA_284), .d1(AA_281), .s2(BB_233_310221), .d2(AA_281), .b(gnd), .g(inst[14]));
NEMR6T g241(.s1(AA_281), .d1(AA_274), .s2(AA_284), .d2(AA_282), .b(gnd), .g(inst[16]));
NEMR6T g242(.s1(AA_274), .d1(AA_242), .s2(AA_340), .d2(AA_451), .b(vdd), .g(inst[13]));
NEMR6T g243(.s1(AA_242), .d1(AA_392), .s2(AA_263), .d2(AA_404), .b(vdd), .g(irq));
NEMR6T g244(.s1(AA_274), .d1(AA_263), .s2(AA_282), .d2(AA_275), .b(gnd), .g(inst[13]));
NEMR6T g245(.s1(AA_263), .d1(AA_262), .s2(AA_275), .d2(AA_264), .b(gnd), .g(irq));
NEMR6T g246(.s1(AA_275), .d1(AA_245), .s2(AA_436), .d2(AA_419), .b(vdd), .g(irq));
NEMR6T g247(.s1(AA_245), .d1(AA_392), .s2(AA_264), .d2(AA_260), .b(gnd), .g(inst[17]));
NEMR6T g248(.s1(stsel[0]), .d1(BB_233_31), .s2(stsel[1]), .d2(BB_286_31), .b(gnd), .g(inst[12]));
NEMR6T g249(.s1(BB_233_31), .d1(BB_233_310), .s2(BB_286_31), .d2(BB_286_310), .b(vdd), .g(z));
NEMR6T g250(.s1(BB_233_310), .d1(AA_285), .s2(BB_233_311), .d2(BB_233_3110), .b(vdd), .g(c));
NEMR6T g251(.s1(AA_285), .d1(AA_283), .s2(BB_233_31011), .d2(AA_253), .b(gnd), .g(inst[10]));
NEMR6T g252(.s1(AA_283), .d1(AA_280), .s2(AA_253), .d2(AA_242), .b(vdd), .g(inst[14]));
NEMR6T g253(.s1(AA_283), .d1(AA_242), .s2(AA_269), .d2(AA_242), .b(vdd), .g(inst[16]));
NEMR6T g254(.s1(AA_283), .d1(AA_282), .s2(AA_269), .d2(AA_282), .b(gnd), .g(inst[16]));
NEMR6T g255(.s1(BB_233_310), .d1(BB_233_3101), .s2(BB_233_311), .d2(BB_233_3111), .b(gnd), .g(c));
NEMR6T g256(.s1(BB_233_3101), .d1(AA_285), .s2(BB_233_3111), .d2(BB_233_31110), .b(vdd), .g(inst[11]));
NEMR6T g257(.s1(BB_233_3101), .d1(BB_233_31011), .s2(BB_233_3110), .d2(BB_233_31101), .b(gnd), .g(inst[11]));
NEMR6T g258(.s1(BB_233_310), .d1(BB_233_310221), .s2(BB_233_31101), .d2(BB_233_311011), .b(gnd), .g(inst[10]));
NEMR6T g259(.s1(BB_233_31), .d1(BB_233_311), .s2(BB_286_31), .d2(BB_286_311), .b(gnd), .g(z));
NEMR6T g260(.s1(BB_233_31101), .d1(AA_242), .s2(BB_233_31120), .d2(AA_283), .b(vdd), .g(inst[10]));
NEMR6T g261(.s1(BB_233_311011), .d1(AA_280), .s2(BB_233_311111), .d2(AA_281), .b(vdd), .g(inst[14]));
NEMR6T g262(.s1(BB_233_3110), .d1(AA_279), .s2(BB_233_31110), .d2(AA_279), .b(gnd), .g(inst[10]));
NEMR6T g263(.s1(AA_279), .d1(AA_269), .s2(BB_233_31120), .d2(AA_281), .b(gnd), .g(inst[14]));
NEMR6T g264(.s1(BB_233_3111), .d1(BB_233_31111), .s2(BB_233_311), .d2(BB_233_31121), .b(gnd), .g(inst[11]));
NEMR6T g265(.s1(BB_233_31111), .d1(BB_233_311111), .s2(BB_233_31120), .d2(AA_253), .b(gnd), .g(inst[10]));
NEMR6T g266(.s1(BB_233_311), .d1(BB_233_31120), .s2(BB_286_3101), .d2(AA_336), .b(vdd), .g(inst[11]));
NEMR6T g267(.s1(BB_233_31121), .d1(BB_233_311211), .s2(BB_233_31211), .d2(AA_279), .b(gnd), .g(inst[10]));
NEMR6T g268(.s1(BB_233_311211), .d1(AA_269), .s2(BB_286_30), .d2(AA_341), .b(vdd), .g(inst[14]));
NEMR6T g269(.s1(BB_233_311211), .d1(AA_281), .s2(BB_286_30), .d2(AA_342), .b(gnd), .g(inst[14]));
NEMR6T g270(.s1(BB_233_31), .d1(BB_233_3121), .s2(BB_286_310), .d2(BB_286_3101), .b(gnd), .g(c));
NEMR6T g271(.s1(BB_233_3121), .d1(BB_233_31211), .s2(BB_286_3101), .d2(BB_286_31011), .b(gnd), .g(inst[11]));
NEMR6T g272(.s1(BB_233_31211), .d1(AA_284), .s2(AA_336), .d2(AA_335), .b(vdd), .g(inst[10]));
NEMR6T g273(.s1(AA_341), .d1(AA_456), .s2(AA_342), .d2(AA_292), .b(vdd), .g(inst[16]));
NEMR6T g274(.s1(AA_456), .d1(AA_436), .s2(AA_341), .d2(AA_461), .b(gnd), .g(inst[13]));
NEMR6T g275(.s1(AA_436), .d1(AA_403), .s2(BB_343_3100), .d2(AA_423), .b(gnd), .g(inst[17]));
NEMR6T g276(.s1(AA_292), .d1(AA_392), .s2(BB_286_30222221), .d2(AA_451), .b(gnd), .g(inst[13]));
NEMR6T g277(.s1(AA_342), .d1(AA_340), .s2(BB_286_30), .d2(BB_286_30222221), .b(gnd), .g(inst[16]));
NEMR6T g278(.s1(BB_286_30), .d1(AA_294), .s2(AA_335), .d2(AA_392), .b(vdd), .g(inst[16]));
NEMR6T g279(.s1(AA_294), .d1(AA_392), .s2(BB_286_30222221), .d2(AA_461), .b(vdd), .g(inst[13]));
NEMR6T g280(.s1(BB_286_310), .d1(AA_336), .s2(BB_286_311), .d2(BB_286_3110), .b(vdd), .g(c));
NEMR6T g281(.s1(AA_335), .d1(AA_334), .s2(AA_325), .d2(AA_341), .b(vdd), .g(inst[14]));
NEMR6T g282(.s1(AA_334), .d1(AA_461), .s2(AA_298), .d2(AA_294), .b(gnd), .g(inst[16]));
NEMR6T g283(.s1(AA_335), .d1(AA_298), .s2(BB_286_310221), .d2(AA_342), .b(gnd), .g(inst[14]));
NEMR6T g284(.s1(AA_336), .d1(AA_325), .s2(BB_286_31011), .d2(AA_326), .b(gnd), .g(inst[10]));
NEMR6T g285(.s1(AA_325), .d1(AA_294), .s2(AA_308), .d2(AA_392), .b(vdd), .g(inst[16]));
NEMR6T g286(.s1(AA_325), .d1(AA_302), .s2(AA_308), .d2(AA_461), .b(gnd), .g(inst[16]));
NEMR6T g287(.s1(AA_302), .d1(AA_461), .s2(BB_286_32222201), .d2(AA_436), .b(vdd), .g(inst[13]));
NEMR6T g288(.s1(AA_326), .d1(AA_308), .s2(BB_286_311011), .d2(AA_341), .b(vdd), .g(inst[14]));
NEMR6T g289(.s1(BB_286_310), .d1(BB_286_310221), .s2(BB_286_31101), .d2(BB_286_311011), .b(gnd), .g(inst[10]));
NEMR6T g290(.s1(BB_286_310), .d1(AA_460), .s2(AA_311), .d2(AA_302), .b(gnd), .g(inst[16]));
NEMR6T g291(.s1(BB_286_3110), .d1(BB_286_31101), .s2(BB_286_3111), .d2(BB_286_31111), .b(gnd), .g(inst[11]));
NEMR6T g292(.s1(BB_286_31101), .d1(AA_335), .s2(BB_286_31111), .d2(AA_313), .b(vdd), .g(inst[10]));
NEMR6T g293(.s1(BB_286_3110), .d1(AA_328), .s2(BB_286_31110), .d2(AA_328), .b(gnd), .g(inst[10]));
NEMR6T g294(.s1(AA_328), .d1(AA_311), .s2(BB_286_311111), .d2(AA_313), .b(gnd), .g(inst[14]));
NEMR6T g295(.s1(AA_311), .d1(AA_294), .s2(BB_286_312110), .d2(AA_294), .b(vdd), .g(inst[16]));
NEMR6T g296(.s1(BB_286_3110), .d1(AA_460), .s2(BB_286_31110), .d2(AA_460), .b(gnd), .g(inst[16]));
NEMR6T g297(.s1(BB_286_311), .d1(BB_286_3111), .s2(BB_286_31), .d2(BB_286_3121), .b(gnd), .g(c));
NEMR6T g298(.s1(BB_286_3111), .d1(BB_286_31110), .s2(BB_286_311), .d2(BB_286_31120), .b(vdd), .g(inst[11]));
NEMR6T g299(.s1(AA_313), .d1(AA_460), .s2(BB_286_312110), .d2(AA_302), .b(gnd), .g(inst[16]));
NEMR6T g300(.s1(BB_286_31111), .d1(BB_286_311111), .s2(BB_286_31120), .d2(AA_326), .b(gnd), .g(inst[10]));
NEMR6T g301(.s1(BB_286_311111), .d1(AA_292), .s2(BB_286_311211), .d2(AA_311), .b(vdd), .g(inst[14]));
NEMR6T g302(.s1(BB_286_31120), .d1(AA_325), .s2(BB_286_31211), .d2(BB_286_312110), .b(vdd), .g(inst[10]));
NEMR6T g303(.s1(BB_286_31120), .d1(AA_342), .s2(BB_286_311211), .d2(AA_342), .b(gnd), .g(inst[14]));
NEMR6T g304(.s1(BB_286_311), .d1(BB_286_31121), .s2(BB_286_3121), .d2(BB_286_31211), .b(gnd), .g(inst[11]));
NEMR6T g305(.s1(BB_286_31121), .d1(BB_286_311211), .s2(BB_286_31211), .d2(AA_328), .b(gnd), .g(inst[10]));
NEMR6T g306(.s1(BB_286_312110), .d1(AA_341), .s2(stsel[1]), .d2(BB_286_3222220), .b(vdd), .g(inst[14]));
NEMR6T g307(.s1(BB_286_312110), .d1(AA_342), .s2(stsel[1]), .d2(BB_286_3222221), .b(gnd), .g(inst[14]));
NEMR6T g308(.s1(BB_286_3222220), .d1(BB_286_32222201), .s2(BB_286_3222221), .d2(BB_286_32222211), .b(gnd), .g(inst[16]));
NEMR6T g309(.s1(BB_286_32222211), .d1(AA_461), .s2(BB_343_311), .d2(AA_453), .b(gnd), .g(inst[13]));
NEMR6T g310(.s1(read_strobe), .d1(AA_392), .s2(write_strobe), .d2(AA_392), .b(vdd), .g(inst[14]));
NEMR6T g311(.s1(read_strobe), .d1(BB_343_31), .s2(BB_350_30), .d2(BB_350_301), .b(gnd), .g(inst[14]));
NEMR6T g312(.s1(BB_343_31), .d1(BB_343_310), .s2(BB_350_301), .d2(BB_350_3010), .b(vdd), .g(inst[16]));
NEMR6T g313(.s1(BB_343_310), .d1(BB_343_3100), .s2(BB_343_311), .d2(AA_392), .b(vdd), .g(inst[13]));
NEMR6T g314(.s1(BB_343_3100), .d1(AA_402), .s2(BB_343_3121), .d2(AA_392), .b(vdd), .g(irq));
NEMR6T g315(.s1(BB_343_310), .d1(AA_420), .s2(BB_343_3121), .d2(BB_343_31211), .b(gnd), .g(irq));
NEMR6T g316(.s1(BB_343_31), .d1(BB_343_311), .s2(BB_350_311), .d2(AA_460), .b(gnd), .g(inst[16]));
NEMR6T g317(.s1(BB_343_31), .d1(BB_343_3121), .s2(BB_350_301), .d2(AA_451), .b(gnd), .g(inst[13]));
NEMR6T g318(.s1(BB_343_31211), .d1(AA_423), .s2(BB_361_301100), .d2(AA_395), .b(gnd), .g(inst[17]));
NEMR4T g319(.s(write_strobe), .d(BB_350_30), .b(vdd), .g(clk));
NEMR6T g320(.s1(BB_350_3010), .d1(AA_436), .s2(BB_361_3011), .d2(BB_361_30110), .b(vdd), .g(inst[13]));
NEMR6T g321(.s1(BB_350_3010), .d1(AA_452), .s2(interrupt_ack), .d2(BB_360_31), .b(gnd), .g(irq));
NEMR4T g322(.s(write_strobe), .d(BB_350_31), .b(gnd), .g(clk));
NEMR6T g323(.s1(BB_350_31), .d1(BB_350_311), .s2(write_strobe), .d2(BB_350_321), .b(gnd), .g(inst[14]));
NEMR6T g324(.s1(BB_350_311), .d1(AA_392), .s2(BB_361_301), .d2(AA_392), .b(vdd), .g(inst[16]));
NEMR6T g325(.s1(BB_350_321), .d1(AA_464), .s2(BB_361_301), .d2(BB_361_3011), .b(gnd), .g(inst[16]));
NEMR6T g326(.s1(interrupt_ack), .d1(AA_392), .s2(BB_361_30110), .d2(BB_361_301100), .b(vdd), .g(irq));
NEMR6T g327(.s1(BB_360_31), .d1(vdd), .s2(AA_372), .d2(AA_394), .b(vdd), .g(ireset));
NEMR6T g328(.s1(BB_360_31), .d1(gnd), .s2(BB_361_312110), .d2(AA_392), .b(gnd), .g(ireset));
NEMR4T g329(.s(next_interrupt_enabled), .d(BB_361_30), .b(vdd), .g(interrupt_enabled));
NEMR6T g330(.s1(BB_361_30), .d1(AA_392), .s2(BB_361_31), .d2(BB_361_310), .b(vdd), .g(inst[0]));
NEMR6T g331(.s1(BB_361_30), .d1(BB_361_301), .s2(BB_361_31), .d2(BB_361_311), .b(gnd), .g(inst[0]));
NEMR6T g332(.s1(BB_361_30110), .d1(AA_392), .s2(BB_361_31010), .d2(AA_422), .b(vdd), .g(inst[17]));
NEMR6T g333(.s1(BB_361_30110), .d1(AA_403), .s2(BB_361_31010), .d2(AA_409), .b(gnd), .g(inst[17]));
NEMR6T g334(.s1(BB_361_3011), .d1(AA_421), .s2(BB_361_3101), .d2(BB_361_31011), .b(gnd), .g(inst[13]));
NEMR6T g335(.s1(BB_361_3011), .d1(AA_452), .s2(BB_361_31010), .d2(AA_401), .b(gnd), .g(irq));
NEMR4T g336(.s(next_interrupt_enabled), .d(BB_361_31), .b(gnd), .g(interrupt_enabled));
NEMR6T g337(.s1(BB_361_310), .d1(BB_361_3101), .s2(BB_361_311), .d2(BB_361_3111), .b(gnd), .g(inst[16]));
NEMR6T g338(.s1(BB_361_3101), .d1(BB_361_31010), .s2(BB_361_3111), .d2(BB_361_31110), .b(vdd), .g(inst[13]));
NEMR6T g339(.s1(BB_361_31010), .d1(AA_434), .s2(BB_361_31110), .d2(AA_422), .b(vdd), .g(irq));
NEMR6T g340(.s1(BB_361_31011), .d1(AA_404), .s2(BB_361_3101), .d2(AA_408), .b(gnd), .g(irq));
NEMR6T g341(.s1(BB_361_31110), .d1(AA_392), .s2(BB_361_3120), .d2(AA_392), .b(gnd), .g(irq));
NEMR6T g342(.s1(BB_361_31), .d1(BB_361_3120), .s2(BB_373_30), .d2(BB_373_300), .b(vdd), .g(inst[16]));
NEMR6T g343(.s1(BB_361_3120), .d1(AA_435), .s2(BB_361_31211), .d2(BB_361_312110), .b(vdd), .g(irq));
NEMR6T g344(.s1(BB_361_31), .d1(BB_361_3121), .s2(BB_361_321), .d2(BB_361_3211), .b(gnd), .g(inst[16]));
NEMR6T g345(.s1(BB_361_3121), .d1(BB_361_31211), .s2(BB_361_3211), .d2(BB_361_32111), .b(gnd), .g(inst[13]));
NEMR6T g346(.s1(BB_361_312110), .d1(AA_372), .s2(BB_361_312120), .d2(BB_361_3121201), .b(gnd), .g(inst[17]));
NEMR6T g347(.s1(BB_361_31211), .d1(AA_452), .s2(BB_361_32111), .d2(AA_407), .b(gnd), .g(irq));
NEMR6T g348(.s1(BB_361_3121), .d1(BB_361_312120), .s2(BB_361_32110), .d2(BB_361_321100), .b(vdd), .g(irq));
NEMR6T g349(.s1(BB_361_312120), .d1(AA_424), .s2(BB_373_31020), .d2(AA_424), .b(vdd), .g(inst[17]));
NEMR6T g350(.s1(BB_361_3121201), .d1(AA_391), .s2(BB_373_30000), .d2(AA_391), .b(vdd), .g(ireset));
NEMR4T g351(.s(next_interrupt_enabled), .d(BB_361_321), .b(gnd), .g(inst[0]));
NEMR6T g352(.s1(BB_361_3211), .d1(BB_361_32110), .s2(BB_373_300), .d2(BB_373_3000), .b(vdd), .g(inst[13]));
NEMR6T g353(.s1(BB_361_321100), .d1(AA_372), .s2(AA_386), .d2(AA_410), .b(gnd), .g(inst[17]));
NEMR6T g354(.s1(werf), .d1(BB_373_30), .s2(wesp), .d2(AA_392), .b(vdd), .g(inst[14]));
NEMR6T g355(.s1(BB_373_3000), .d1(BB_373_30000), .s2(AA_386), .d2(AA_406), .b(vdd), .g(irq));
NEMR6T g356(.s1(BB_373_30000), .d1(AA_395), .s2(BB_373_31020), .d2(AA_392), .b(gnd), .g(ireset));
NEMR4T g357(.s(BB_373_30000), .d(gnd), .b(gnd), .g(inst[15]));
NEMR6T g358(.s1(BB_373_3000), .d1(AA_392), .s2(AA_386), .d2(AA_407), .b(gnd), .g(irq));
NEMR6T g359(.s1(BB_373_30), .d1(AA_386), .s2(BB_373_311), .d2(AA_386), .b(gnd), .g(inst[13]));
NEMR6T g360(.s1(werf), .d1(BB_373_31), .s2(wesp), .d2(BB_387_31), .b(gnd), .g(inst[14]));
NEMR6T g361(.s1(BB_373_31), .d1(BB_373_310), .s2(BB_387_31), .d2(AA_456), .b(vdd), .g(inst[16]));
NEMR4T g362(.s(BB_373_310), .d(BB_373_31020), .b(vdd), .g(irq));
NEMR4T g363(.s(BB_373_310), .d(AA_454), .b(gnd), .g(irq));
NEMR4T g364(.s(BB_373_310), .d(AA_401), .b(gnd), .g(inst[17]));
NEMR6T g365(.s1(BB_373_31), .d1(BB_373_311), .s2(werf), .d2(BB_373_321), .b(gnd), .g(inst[16]));
NEMR6T g366(.s1(BB_373_321), .d1(AA_386), .s2(BB_387_31), .d2(AA_392), .b(vdd), .g(inst[13]));
NEMR4T g367(.s(BB_387_31), .d(AA_460), .b(gnd), .g(inst[16]));
NEMR4T g368(.s(BB_387_31), .d(AA_461), .b(gnd), .g(inst[13]));
