module Instruction_decode(clk, ireset, irq, inst, c, z, read_strobe,
     write_strobe, interrupt_ack, next_interrupt_enabled,
     interrupt_enabled, zsel, csel, wsel, pcsel, stsel, werf, wesp);
  input clk, ireset, irq, c, z, interrupt_enabled;
  input [17:0] inst;
  output read_strobe, write_strobe, interrupt_ack,
       next_interrupt_enabled, werf, wesp;
  output [2:0] zsel, csel, wsel;
  output [1:0] pcsel, stsel;


  wire csel[0], csel[0]0, csel[0]00, csel[0]000, csel[0]01, csel[0]011, csel[0]1, csel[0]10, csel[0]100, csel[0]1000, 
  csel[0]10000, csel[0]100001, csel[0]11, csel[0]120, csel[0]20, csel[0]200, csel[0]2000, csel[0]21, csel[0]210, csel[0]2100, 
  csel[0]21000, csel[0]220, csel[0]2201, csel[0]22010, csel[0]220100, csel[0]220101, csel[0]221, csel[0]22120, csel[0]221200, csel[1], 
  csel[1]0, csel[1]00, csel[1]000, csel[1]0000, csel[1]00000, csel[1]1, csel[1]10, csel[1]100, csel[1]1000, csel[1]20, 
  csel[1]200, csel[1]2000, csel[1]20000, csel[1]201, csel[1]2010, csel[1]20100, csel[1]2011, csel[1]21, csel[1]210, csel[1]2100, 
  csel[1]21001, csel[1]2120, csel[1]21200, csel[1]221, csel[1]2210, csel[1]22101, csel[1]2221, csel[2], csel[2]0, csel[2]00, 
  csel[2]000, csel[2]0000, csel[2]00000, csel[2]001, csel[2]0010, csel[2]00100, csel[2]01, csel[2]011, csel[2]0110, csel[2]01100, 
  csel[2]0120, csel[2]1, csel[2]120, csel[2]121, csel[2]220, csel[2]2200, int_0, int_1, int_101, int_102, 
  int_103, int_104, int_105, int_107, int_108, int_109, int_11, int_110, int_112, int_113, 
  int_114, int_115, int_116, int_117, int_118, int_12, int_120, int_121, int_122, int_123, 
  int_124, int_126, int_127, int_128, int_129, int_13, int_130, int_131, int_132, int_133, 
  int_134, int_135, int_136, int_139, int_140, int_141, int_143, int_144, int_145, int_146, 
  int_147, int_148, int_149, int_15, int_150, int_151, int_152, int_153, int_154, int_155, 
  int_156, int_157, int_158, int_159, int_16, int_160, int_162, int_163, int_164, int_165, 
  int_166, int_167, int_168, int_171, int_172, int_173, int_174, int_175, int_176, int_177, 
  int_178, int_179, int_180, int_181, int_182, int_183, int_184, int_185, int_186, int_187, 
  int_188, int_189, int_19, int_190, int_191, int_192, int_193, int_194, int_195, int_196, 
  int_197, int_198, int_199, int_2, int_20, int_200, int_201, int_202, int_203, int_204, 
  int_205, int_206, int_207, int_208, int_209, int_21, int_210, int_211, int_212, int_213, 
  int_214, int_215, int_216, int_217, int_218, int_219, int_22, int_220, int_221, int_222, 
  int_223, int_224, int_225, int_226, int_24, int_25, int_26, int_27, int_29, int_3, 
  int_31, int_32, int_33, int_34, int_35, int_36, int_37, int_38, int_39, int_4, 
  int_40, int_41, int_42, int_43, int_49, int_50, int_51, int_52, int_55, int_56, 
  int_58, int_59, int_6, int_60, int_61, int_62, int_63, int_64, int_66, int_67, 
  int_68, int_69, int_70, int_71, int_72, int_73, int_75, int_78, int_8, int_82, 
  int_84, int_86, int_87, int_88, int_89, int_9, int_90, int_91, int_92, int_93, 
  int_94, int_97, int_98, int_99, next_interrupt_enabled, next_interrupt_enabled0, next_interrupt_enabled00, next_interrupt_enabled001, next_interrupt_enabled1, next_interrupt_enabled10, 
  next_interrupt_enabled12220, next_interrupt_enabled122200, next_interrupt_enabled20, next_interrupt_enabled201, pcsel[0], pcsel[0]0, pcsel[0]00, pcsel[0]000, pcsel[0]001, pcsel[0]01, 
  pcsel[0]010, pcsel[0]021, pcsel[0]1, pcsel[0]10, pcsel[0]100, pcsel[0]101, pcsel[0]11, pcsel[0]110, pcsel[0]121, pcsel[0]20, 
  pcsel[0]200, pcsel[0]21, pcsel[0]221, pcsel[1], pcsel[1]0, pcsel[1]00, pcsel[1]000, pcsel[1]001, pcsel[1]01, pcsel[1]010, 
  pcsel[1]021, pcsel[1]1, pcsel[1]10, pcsel[1]100, pcsel[1]101, pcsel[1]11, pcsel[1]110, pcsel[1]121, pcsel[1]20, pcsel[1]200, 
  pcsel[1]21, pcsel[1]221, read_strobe, read_strobe0, read_strobe00, read_strobe000, read_strobe0000, read_strobe00000, read_strobe01, read_strobe1, 
  stsel[0], stsel[0]0, stsel[0]00, stsel[0]000, stsel[0]001, stsel[0]01, stsel[0]010, stsel[0]021, stsel[0]1, stsel[0]10, 
  stsel[0]100, stsel[0]10020, stsel[0]101, stsel[0]11, stsel[0]110, stsel[0]121, stsel[0]20, stsel[0]200, stsel[0]200220, stsel[0]201, 
  stsel[0]21, stsel[0]210, stsel[0]221, stsel[1], stsel[1]0, stsel[1]00, stsel[1]000, stsel[1]001, stsel[1]01, stsel[1]010, 
  stsel[1]021, stsel[1]1, stsel[1]10, stsel[1]100, stsel[1]10020, stsel[1]100200, stsel[1]101, stsel[1]11, stsel[1]110, stsel[1]121, 
  stsel[1]20, stsel[1]200, stsel[1]200220, stsel[1]2002200, stsel[1]21, stsel[1]221, werf, werf0, werf00, werf000, 
  werf0001, werf00010, werf01, werf011, werf021, werf1, werf10, werf100, werf1000, werf11, 
  werf20, werf200, werf2000, werf20000, werf200000, werf20001, wesp, wesp0, wesp00, wesp001, 
  wesp0011, wesp00110, wesp001101, wesp01, wesp011, wesp021, wesp1, write_strobe, write_strobe0, write_strobe00, 
  write_strobe000, write_strobe0000, write_strobe00000, write_strobe000001, write_strobe1, write_strobe10, write_strobe101, write_strobe11, write_strobe20, wsel[0], 
  wsel[0]0, wsel[0]01, wsel[1], wsel[1]0, zsel[0], zsel[0]0, zsel[0]00, zsel[0]000, zsel[0]0000, zsel[0]001, 
  zsel[0]0011, zsel[0]01, zsel[0]011, zsel[0]1, zsel[0]121, zsel[0]1210, zsel[0]1211, zsel[0]12120, zsel[0]1220, zsel[0]220, 
  zsel[1], zsel[1]0, zsel[1]00, zsel[1]000, zsel[1]0000, zsel[1]00000, zsel[1]0020, zsel[1]01, zsel[1]010, zsel[1]0100, 
  zsel[1]0101, zsel[1]011, zsel[1]0110, zsel[1]1, zsel[1]120, zsel[1]121, zsel[1]1210, zsel[1]1220, zsel[1]220, zsel[1]2200, 
  zsel[1]221, zsel[1]2211, zsel[1]2220, zsel[2], zsel[2]0, zsel[2]00, zsel[2]000, zsel[2]1, zsel[2]10, zsel[2]101, 
  zsel[2]11, zsel[2]20;


  assign wsel[2] = inst[16];

NEMR4T g1(.s(zsel[0]), .d(zsel[0]0), .b(vdd), .g(inst[13]));
NEMR4T g2(.s(zsel[0]0), .d(zsel[0]00), .b(vdd), .g(inst[14]));
NEMR4T g3(.s(zsel[0]00), .d(zsel[0]000), .b(vdd), .g(inst[16]));
NEMR4T g4(.s(zsel[0]000), .d(zsel[0]0000), .b(vdd), .g(inst[15]));
NEMR4T g5(.s(zsel[0]0000), .d(int_139), .b(vdd), .g(irq));
NEMR4T g6(.s(int_139), .d(int_0), .b(gnd), .g(inst[17]));
NEMR4T g7(.s(int_0), .d(vdd), .b(gnd), .g(vdd));
NEMR4T g8(.s(zsel[0]00), .d(zsel[0]001), .b(gnd), .g(inst[16]));
NEMR4T g9(.s(zsel[0]001), .d(int_1), .b(vdd), .g(inst[15]));
NEMR4T g10(.s(int_1), .d(gnd), .b(vdd), .g(ireset));
NEMR4T g11(.s(zsel[0]001), .d(zsel[0]0011), .b(gnd), .g(inst[15]));
NEMR4T g12(.s(zsel[0]0011), .d(int_140), .b(vdd), .g(irq));
NEMR4T g13(.s(int_140), .d(int_2), .b(vdd), .g(inst[17]));
NEMR4T g14(.s(int_2), .d(vdd), .b(vdd), .g(ireset));
NEMR4T g15(.s(zsel[0]0011), .d(int_3), .b(gnd), .g(irq));
NEMR4T g16(.s(int_3), .d(int_1), .b(vdd), .g(inst[17]));
NEMR4T g17(.s(zsel[0]0011), .d(int_1), .b(gnd), .g(inst[17]));
NEMR4T g18(.s(zsel[0]001), .d(vdd), .b(gnd), .g(ireset));
NEMR4T g19(.s(zsel[0]0), .d(zsel[0]01), .b(gnd), .g(inst[14]));
NEMR4T g20(.s(zsel[0]01), .d(zsel[0]011), .b(gnd), .g(inst[16]));
NEMR4T g21(.s(zsel[0]011), .d(int_198), .b(vdd), .g(inst[15]));
NEMR4T g22(.s(int_198), .d(int_141), .b(gnd), .g(irq));
NEMR4T g23(.s(int_141), .d(int_4), .b(gnd), .g(inst[17]));
NEMR4T g24(.s(int_4), .d(gnd), .b(vdd), .g(ireset));
NEMR4T g25(.s(int_4), .d(vdd), .b(gnd), .g(ireset));
NEMR4T g26(.s(zsel[0]011), .d(int_140), .b(vdd), .g(irq));
NEMR4T g27(.s(zsel[0]011), .d(int_3), .b(gnd), .g(irq));
NEMR4T g28(.s(zsel[0]011), .d(int_6), .b(vdd), .g(inst[17]));
NEMR4T g29(.s(int_6), .d(vdd), .b(gnd), .g(ireset));
NEMR4T g30(.s(zsel[0]01), .d(int_198), .b(gnd), .g(inst[15]));
NEMR4T g31(.s(zsel[0]01), .d(int_141), .b(vdd), .g(irq));
NEMR4T g32(.s(zsel[0]), .d(zsel[0]1), .b(gnd), .g(inst[13]));
NEMR4T g33(.s(zsel[0]1), .d(int_143), .b(gnd), .g(inst[14]));
NEMR4T g34(.s(int_143), .d(int_8), .b(vdd), .g(inst[16]));
NEMR4T g35(.s(int_8), .d(int_141), .b(gnd), .g(inst[15]));
NEMR4T g36(.s(zsel[0]1), .d(zsel[0]121), .b(gnd), .g(inst[16]));
NEMR4T g37(.s(zsel[0]121), .d(zsel[0]1210), .b(vdd), .g(inst[15]));
NEMR4T g38(.s(zsel[0]1210), .d(int_3), .b(vdd), .g(irq));
NEMR4T g39(.s(zsel[0]1210), .d(int_4), .b(gnd), .g(irq));
NEMR4T g40(.s(zsel[0]121), .d(zsel[0]1211), .b(gnd), .g(inst[15]));
NEMR4T g41(.s(zsel[0]1211), .d(int_140), .b(vdd), .g(irq));
NEMR4T g42(.s(zsel[0]1211), .d(int_9), .b(gnd), .g(irq));
NEMR4T g43(.s(int_9), .d(int_4), .b(vdd), .g(inst[17]));
NEMR4T g44(.s(zsel[0]1211), .d(int_4), .b(gnd), .g(inst[17]));
NEMR4T g45(.s(zsel[0]121), .d(zsel[0]12120), .b(vdd), .g(irq));
NEMR4T g46(.s(zsel[0]12120), .d(int_6), .b(vdd), .g(inst[17]));
NEMR4T g47(.s(zsel[0]1), .d(zsel[0]1220), .b(vdd), .g(inst[15]));
NEMR4T g48(.s(zsel[0]1220), .d(int_141), .b(vdd), .g(irq));
NEMR4T g49(.s(zsel[0]), .d(int_143), .b(vdd), .g(inst[14]));
NEMR4T g50(.s(zsel[0]), .d(zsel[0]220), .b(vdd), .g(inst[16]));
NEMR4T g51(.s(zsel[0]220), .d(int_198), .b(vdd), .g(inst[15]));
NEMR4T g52(.s(zsel[0]220), .d(int_4), .b(vdd), .g(inst[17]));
NEMR4T g53(.s(zsel[1]), .d(zsel[1]0), .b(vdd), .g(inst[14]));
NEMR4T g54(.s(zsel[1]0), .d(zsel[1]00), .b(vdd), .g(inst[13]));
NEMR4T g55(.s(zsel[1]00), .d(zsel[1]000), .b(vdd), .g(inst[15]));
NEMR4T g56(.s(zsel[1]000), .d(zsel[1]0000), .b(vdd), .g(inst[16]));
NEMR4T g57(.s(zsel[1]0000), .d(zsel[1]00000), .b(vdd), .g(irq));
NEMR4T g58(.s(zsel[1]00000), .d(int_11), .b(vdd), .g(ireset));
NEMR4T g59(.s(int_11), .d(vdd), .b(gnd), .g(inst[17]));
NEMR4T g60(.s(zsel[1]00), .d(zsel[1]0020), .b(vdd), .g(inst[16]));
NEMR4T g61(.s(zsel[1]0020), .d(int_144), .b(vdd), .g(irq));
NEMR4T g62(.s(int_144), .d(int_12), .b(vdd), .g(ireset));
NEMR4T g63(.s(int_12), .d(gnd), .b(vdd), .g(inst[17]));
NEMR4T g64(.s(zsel[1]0020), .d(int_145), .b(gnd), .g(irq));
NEMR4T g65(.s(int_145), .d(int_13), .b(vdd), .g(ireset));
NEMR4T g66(.s(int_13), .d(gnd), .b(gnd), .g(vdd));
NEMR4T g67(.s(zsel[1]0020), .d(int_12), .b(gnd), .g(ireset));
NEMR4T g68(.s(zsel[1]0), .d(zsel[1]01), .b(gnd), .g(inst[13]));
NEMR4T g69(.s(zsel[1]01), .d(zsel[1]010), .b(vdd), .g(inst[15]));
NEMR4T g70(.s(zsel[1]010), .d(zsel[1]0100), .b(vdd), .g(inst[16]));
NEMR4T g71(.s(zsel[1]0100), .d(int_144), .b(vdd), .g(irq));
NEMR4T g72(.s(zsel[1]010), .d(zsel[1]0101), .b(gnd), .g(inst[16]));
NEMR4T g73(.s(zsel[1]0101), .d(int_146), .b(vdd), .g(irq));
NEMR4T g74(.s(int_146), .d(int_15), .b(vdd), .g(ireset));
NEMR4T g75(.s(int_15), .d(vdd), .b(vdd), .g(inst[17]));
NEMR4T g76(.s(zsel[1]0101), .d(int_16), .b(gnd), .g(ireset));
NEMR4T g77(.s(int_16), .d(gnd), .b(gnd), .g(inst[17]));
NEMR4T g78(.s(zsel[1]010), .d(int_144), .b(gnd), .g(irq));
NEMR4T g79(.s(zsel[1]010), .d(int_16), .b(vdd), .g(ireset));
NEMR4T g80(.s(zsel[1]010), .d(int_12), .b(gnd), .g(ireset));
NEMR4T g81(.s(zsel[1]01), .d(zsel[1]011), .b(gnd), .g(inst[15]));
NEMR4T g82(.s(zsel[1]011), .d(zsel[1]0110), .b(vdd), .g(inst[16]));
NEMR4T g83(.s(zsel[1]0110), .d(int_146), .b(vdd), .g(irq));
NEMR4T g84(.s(zsel[1]0110), .d(int_145), .b(gnd), .g(irq));
NEMR4T g85(.s(zsel[1]0110), .d(int_12), .b(gnd), .g(ireset));
NEMR4T g86(.s(zsel[1]), .d(zsel[1]1), .b(gnd), .g(inst[14]));
NEMR4T g87(.s(zsel[1]1), .d(int_199), .b(gnd), .g(inst[13]));
NEMR4T g88(.s(int_199), .d(int_147), .b(vdd), .g(inst[15]));
NEMR4T g89(.s(int_147), .d(int_21), .b(gnd), .g(inst[16]));
NEMR4T g90(.s(int_21), .d(int_19), .b(vdd), .g(irq));
NEMR4T g91(.s(int_19), .d(int_12), .b(vdd), .g(ireset));
NEMR4T g92(.s(int_19), .d(gnd), .b(gnd), .g(inst[17]));
NEMR4T g93(.s(int_21), .d(int_20), .b(gnd), .g(irq));
NEMR4T g94(.s(int_20), .d(int_13), .b(vdd), .g(ireset));
NEMR4T g95(.s(int_20), .d(int_16), .b(gnd), .g(ireset));
NEMR4T g96(.s(int_21), .d(int_12), .b(gnd), .g(ireset));
NEMR4T g97(.s(zsel[1]1), .d(zsel[1]120), .b(vdd), .g(inst[15]));
NEMR4T g98(.s(zsel[1]120), .d(int_145), .b(vdd), .g(inst[16]));
NEMR4T g99(.s(zsel[1]1), .d(zsel[1]121), .b(gnd), .g(inst[15]));
NEMR4T g100(.s(zsel[1]121), .d(zsel[1]1210), .b(vdd), .g(inst[16]));
NEMR4T g101(.s(zsel[1]1210), .d(int_146), .b(vdd), .g(irq));
NEMR4T g102(.s(zsel[1]1210), .d(int_145), .b(gnd), .g(irq));
NEMR4T g103(.s(zsel[1]1), .d(zsel[1]1220), .b(vdd), .g(inst[16]));
NEMR4T g104(.s(zsel[1]1220), .d(int_12), .b(gnd), .g(ireset));
NEMR4T g105(.s(zsel[1]), .d(int_199), .b(vdd), .g(inst[13]));
NEMR4T g106(.s(zsel[1]), .d(zsel[1]220), .b(vdd), .g(inst[15]));
NEMR4T g107(.s(zsel[1]220), .d(zsel[1]2200), .b(vdd), .g(inst[16]));
NEMR4T g108(.s(zsel[1]2200), .d(int_22), .b(vdd), .g(irq));
NEMR4T g109(.s(int_22), .d(int_16), .b(gnd), .g(ireset));
NEMR4T g110(.s(zsel[1]), .d(zsel[1]221), .b(gnd), .g(inst[15]));
NEMR4T g111(.s(zsel[1]221), .d(zsel[1]2211), .b(gnd), .g(inst[16]));
NEMR4T g112(.s(zsel[1]2211), .d(int_144), .b(vdd), .g(irq));
NEMR4T g113(.s(zsel[1]2211), .d(int_20), .b(gnd), .g(irq));
NEMR4T g114(.s(zsel[1]2211), .d(int_12), .b(gnd), .g(ireset));
NEMR4T g115(.s(zsel[1]221), .d(int_16), .b(vdd), .g(irq));
NEMR4T g116(.s(zsel[1]), .d(zsel[1]2220), .b(vdd), .g(inst[16]));
NEMR4T g117(.s(zsel[1]2220), .d(int_22), .b(gnd), .g(irq));
NEMR4T g118(.s(zsel[2]), .d(zsel[2]0), .b(vdd), .g(inst[14]));
NEMR4T g119(.s(zsel[2]0), .d(zsel[2]00), .b(vdd), .g(inst[13]));
NEMR4T g120(.s(zsel[2]00), .d(zsel[2]000), .b(vdd), .g(irq));
NEMR4T g121(.s(zsel[2]000), .d(int_4), .b(vdd), .g(inst[16]));
NEMR4T g122(.s(zsel[2]000), .d(int_148), .b(gnd), .g(inst[16]));
NEMR4T g123(.s(int_148), .d(int_4), .b(vdd), .g(inst[15]));
NEMR4T g124(.s(int_148), .d(int_139), .b(gnd), .g(inst[15]));
NEMR4T g125(.s(zsel[2]0), .d(int_25), .b(gnd), .g(inst[13]));
NEMR4T g126(.s(int_25), .d(int_24), .b(vdd), .g(inst[16]));
NEMR4T g127(.s(int_24), .d(int_9), .b(gnd), .g(inst[15]));
NEMR4T g128(.s(int_25), .d(int_9), .b(vdd), .g(inst[15]));
NEMR4T g129(.s(int_25), .d(int_4), .b(gnd), .g(inst[17]));
NEMR4T g130(.s(zsel[2]0), .d(int_24), .b(gnd), .g(inst[16]));
NEMR4T g131(.s(zsel[2]), .d(zsel[2]1), .b(gnd), .g(inst[14]));
NEMR4T g132(.s(zsel[2]1), .d(zsel[2]10), .b(vdd), .g(inst[13]));
NEMR4T g133(.s(zsel[2]10), .d(zsel[2]101), .b(gnd), .g(irq));
NEMR4T g134(.s(zsel[2]101), .d(int_24), .b(gnd), .g(inst[16]));
NEMR4T g135(.s(zsel[2]1), .d(zsel[2]11), .b(gnd), .g(inst[13]));
NEMR4T g136(.s(zsel[2]11), .d(int_4), .b(gnd), .g(irq));
NEMR4T g137(.s(zsel[2]1), .d(int_4), .b(vdd), .g(irq));
NEMR4T g138(.s(zsel[2]), .d(zsel[2]20), .b(vdd), .g(inst[13]));
NEMR4T g139(.s(zsel[2]20), .d(int_25), .b(gnd), .g(irq));
NEMR4T g140(.s(csel[0]), .d(csel[0]0), .b(vdd), .g(inst[3]));
NEMR4T g141(.s(csel[0]0), .d(csel[0]00), .b(vdd), .g(inst[16]));
NEMR4T g142(.s(csel[0]00), .d(csel[0]000), .b(vdd), .g(inst[14]));
NEMR4T g143(.s(csel[0]000), .d(int_149), .b(vdd), .g(inst[13]));
NEMR4T g144(.s(int_149), .d(int_26), .b(gnd), .g(inst[17]));
NEMR4T g145(.s(int_26), .d(int_4), .b(vdd), .g(inst[15]));
NEMR4T g146(.s(csel[0]0), .d(csel[0]01), .b(gnd), .g(inst[16]));
NEMR4T g147(.s(csel[0]01), .d(csel[0]011), .b(gnd), .g(inst[14]));
NEMR4T g148(.s(csel[0]011), .d(int_200), .b(vdd), .g(inst[13]));
NEMR4T g149(.s(int_200), .d(int_150), .b(gnd), .g(irq));
NEMR4T g150(.s(int_150), .d(int_27), .b(gnd), .g(inst[17]));
NEMR4T g151(.s(int_27), .d(int_4), .b(gnd), .g(inst[15]));
NEMR4T g152(.s(csel[0]01), .d(int_151), .b(vdd), .g(inst[13]));
NEMR4T g153(.s(int_151), .d(int_149), .b(gnd), .g(irq));
NEMR4T g154(.s(csel[0]), .d(csel[0]1), .b(gnd), .g(inst[3]));
NEMR4T g155(.s(csel[0]1), .d(csel[0]10), .b(vdd), .g(inst[16]));
NEMR4T g156(.s(csel[0]10), .d(csel[0]100), .b(vdd), .g(inst[14]));
NEMR4T g157(.s(csel[0]100), .d(csel[0]1000), .b(vdd), .g(inst[13]));
NEMR4T g158(.s(csel[0]1000), .d(csel[0]10000), .b(vdd), .g(irq));
NEMR4T g159(.s(csel[0]10000), .d(csel[0]100001), .b(gnd), .g(inst[17]));
NEMR4T g160(.s(csel[0]100001), .d(int_0), .b(vdd), .g(inst[15]));
NEMR4T g161(.s(csel[0]1), .d(csel[0]11), .b(gnd), .g(inst[16]));
NEMR4T g162(.s(csel[0]11), .d(int_29), .b(gnd), .g(inst[14]));
NEMR4T g163(.s(int_29), .d(int_198), .b(vdd), .g(inst[13]));
NEMR4T g164(.s(csel[0]1), .d(csel[0]120), .b(vdd), .g(inst[14]));
NEMR4T g165(.s(csel[0]120), .d(int_151), .b(vdd), .g(inst[13]));
NEMR4T g166(.s(csel[0]), .d(csel[0]20), .b(vdd), .g(inst[16]));
NEMR4T g167(.s(csel[0]20), .d(csel[0]200), .b(vdd), .g(inst[14]));
NEMR4T g168(.s(csel[0]200), .d(csel[0]2000), .b(vdd), .g(inst[13]));
NEMR4T g169(.s(csel[0]2000), .d(int_9), .b(vdd), .g(irq));
NEMR4T g170(.s(csel[0]2000), .d(int_27), .b(gnd), .g(inst[17]));
NEMR4T g171(.s(csel[0]200), .d(int_200), .b(gnd), .g(inst[13]));
NEMR4T g172(.s(csel[0]20), .d(int_29), .b(gnd), .g(inst[14]));
NEMR4T g173(.s(csel[0]), .d(csel[0]21), .b(gnd), .g(inst[16]));
NEMR4T g174(.s(csel[0]21), .d(csel[0]210), .b(vdd), .g(inst[14]));
NEMR4T g175(.s(csel[0]210), .d(csel[0]2100), .b(vdd), .g(inst[13]));
NEMR4T g176(.s(csel[0]2100), .d(csel[0]21000), .b(vdd), .g(irq));
NEMR4T g177(.s(csel[0]21000), .d(int_1), .b(vdd), .g(inst[15]));
NEMR4T g178(.s(csel[0]21000), .d(int_2), .b(gnd), .g(inst[15]));
NEMR4T g179(.s(csel[0]21000), .d(vdd), .b(gnd), .g(ireset));
NEMR4T g180(.s(csel[0]210), .d(int_150), .b(gnd), .g(irq));
NEMR4T g181(.s(csel[0]), .d(csel[0]220), .b(vdd), .g(inst[14]));
NEMR4T g182(.s(csel[0]220), .d(csel[0]2201), .b(gnd), .g(inst[13]));
NEMR4T g183(.s(csel[0]2201), .d(csel[0]22010), .b(vdd), .g(irq));
NEMR4T g184(.s(csel[0]22010), .d(csel[0]220100), .b(vdd), .g(inst[17]));
NEMR4T g185(.s(csel[0]220100), .d(int_4), .b(vdd), .g(inst[15]));
NEMR4T g186(.s(csel[0]220100), .d(int_2), .b(gnd), .g(inst[15]));
NEMR4T g187(.s(csel[0]22010), .d(csel[0]220101), .b(gnd), .g(inst[17]));
NEMR4T g188(.s(csel[0]220101), .d(int_1), .b(gnd), .g(inst[15]));
NEMR4T g189(.s(csel[0]22010), .d(int_6), .b(gnd), .g(inst[15]));
NEMR4T g190(.s(csel[0]2201), .d(int_26), .b(gnd), .g(inst[17]));
NEMR4T g191(.s(csel[0]), .d(csel[0]221), .b(gnd), .g(inst[14]));
NEMR4T g192(.s(csel[0]221), .d(int_198), .b(gnd), .g(inst[13]));
NEMR4T g193(.s(csel[0]221), .d(csel[0]22120), .b(vdd), .g(irq));
NEMR4T g194(.s(csel[0]22120), .d(csel[0]221200), .b(vdd), .g(inst[17]));
NEMR4T g195(.s(csel[0]221200), .d(int_1), .b(vdd), .g(inst[15]));
NEMR4T g196(.s(csel[0]221200), .d(int_2), .b(gnd), .g(inst[15]));
NEMR4T g197(.s(csel[0]22120), .d(int_1), .b(gnd), .g(inst[17]));
NEMR4T g198(.s(csel[0]22120), .d(vdd), .b(gnd), .g(ireset));
NEMR4T g199(.s(csel[0]), .d(int_9), .b(gnd), .g(irq));
NEMR4T g200(.s(csel[1]), .d(csel[1]0), .b(vdd), .g(inst[3]));
NEMR4T g201(.s(csel[1]0), .d(csel[1]00), .b(vdd), .g(inst[14]));
NEMR4T g202(.s(csel[1]00), .d(csel[1]000), .b(vdd), .g(inst[13]));
NEMR4T g203(.s(csel[1]000), .d(csel[1]0000), .b(vdd), .g(irq));
NEMR4T g204(.s(csel[1]0000), .d(csel[1]00000), .b(vdd), .g(inst[16]));
NEMR4T g205(.s(csel[1]00000), .d(int_139), .b(vdd), .g(inst[15]));
NEMR4T g206(.s(csel[1]), .d(csel[1]1), .b(gnd), .g(inst[3]));
NEMR4T g207(.s(csel[1]1), .d(csel[1]10), .b(vdd), .g(inst[14]));
NEMR4T g208(.s(csel[1]10), .d(csel[1]100), .b(vdd), .g(inst[13]));
NEMR4T g209(.s(csel[1]100), .d(csel[1]1000), .b(vdd), .g(irq));
NEMR4T g210(.s(csel[1]1000), .d(int_31), .b(vdd), .g(inst[16]));
NEMR4T g211(.s(int_31), .d(int_141), .b(vdd), .g(inst[15]));
NEMR4T g212(.s(csel[1]), .d(csel[1]20), .b(vdd), .g(inst[14]));
NEMR4T g213(.s(csel[1]20), .d(csel[1]200), .b(vdd), .g(inst[13]));
NEMR4T g214(.s(csel[1]200), .d(csel[1]2000), .b(vdd), .g(irq));
NEMR4T g215(.s(csel[1]2000), .d(csel[1]20000), .b(vdd), .g(inst[16]));
NEMR4T g216(.s(csel[1]20000), .d(int_9), .b(vdd), .g(inst[15]));
NEMR4T g217(.s(csel[1]20000), .d(int_4), .b(gnd), .g(inst[15]));
NEMR4T g218(.s(csel[1]2000), .d(int_148), .b(gnd), .g(inst[16]));
NEMR4T g219(.s(csel[1]20), .d(csel[1]201), .b(gnd), .g(inst[13]));
NEMR4T g220(.s(csel[1]201), .d(csel[1]2010), .b(vdd), .g(irq));
NEMR4T g221(.s(csel[1]2010), .d(csel[1]20100), .b(vdd), .g(inst[16]));
NEMR4T g222(.s(csel[1]20100), .d(int_32), .b(gnd), .g(inst[15]));
NEMR4T g223(.s(int_32), .d(int_0), .b(vdd), .g(inst[17]));
NEMR4T g224(.s(csel[1]2010), .d(int_31), .b(gnd), .g(inst[16]));
NEMR4T g225(.s(csel[1]201), .d(csel[1]2011), .b(gnd), .g(irq));
NEMR4T g226(.s(csel[1]2011), .d(int_26), .b(gnd), .g(inst[16]));
NEMR4T g227(.s(csel[1]201), .d(int_26), .b(vdd), .g(inst[16]));
NEMR4T g228(.s(csel[1]201), .d(int_141), .b(gnd), .g(inst[15]));
NEMR4T g229(.s(csel[1]), .d(csel[1]21), .b(gnd), .g(inst[14]));
NEMR4T g230(.s(csel[1]21), .d(csel[1]210), .b(vdd), .g(inst[13]));
NEMR4T g231(.s(csel[1]210), .d(csel[1]2100), .b(vdd), .g(irq));
NEMR4T g232(.s(csel[1]2100), .d(csel[1]21001), .b(gnd), .g(inst[16]));
NEMR4T g233(.s(csel[1]21001), .d(int_32), .b(vdd), .g(inst[15]));
NEMR4T g234(.s(csel[1]21), .d(int_152), .b(gnd), .g(inst[13]));
NEMR4T g235(.s(int_152), .d(int_33), .b(gnd), .g(irq));
NEMR4T g236(.s(int_33), .d(int_9), .b(vdd), .g(inst[15]));
NEMR4T g237(.s(int_33), .d(int_4), .b(gnd), .g(inst[17]));
NEMR4T g238(.s(csel[1]21), .d(csel[1]2120), .b(vdd), .g(irq));
NEMR4T g239(.s(csel[1]2120), .d(csel[1]21200), .b(vdd), .g(inst[16]));
NEMR4T g240(.s(csel[1]21200), .d(int_4), .b(vdd), .g(inst[15]));
NEMR4T g241(.s(csel[1]21200), .d(int_32), .b(gnd), .g(inst[15]));
NEMR4T g242(.s(csel[1]2120), .d(int_31), .b(gnd), .g(inst[16]));
NEMR4T g243(.s(csel[1]2120), .d(int_141), .b(gnd), .g(inst[15]));
NEMR4T g244(.s(csel[1]), .d(int_152), .b(vdd), .g(inst[13]));
NEMR4T g245(.s(csel[1]), .d(csel[1]221), .b(gnd), .g(inst[13]));
NEMR4T g246(.s(csel[1]221), .d(csel[1]2210), .b(vdd), .g(irq));
NEMR4T g247(.s(csel[1]2210), .d(csel[1]22101), .b(gnd), .g(inst[16]));
NEMR4T g248(.s(csel[1]22101), .d(int_9), .b(vdd), .g(inst[15]));
NEMR4T g249(.s(csel[1]), .d(csel[1]2221), .b(gnd), .g(irq));
NEMR4T g250(.s(csel[1]2221), .d(int_24), .b(vdd), .g(inst[16]));
NEMR4T g251(.s(csel[1]), .d(int_24), .b(gnd), .g(inst[16]));
NEMR4T g252(.s(csel[2]), .d(csel[2]0), .b(vdd), .g(inst[14]));
NEMR4T g253(.s(csel[2]0), .d(csel[2]00), .b(vdd), .g(inst[13]));
NEMR4T g254(.s(csel[2]00), .d(csel[2]000), .b(vdd), .g(inst[16]));
NEMR4T g255(.s(csel[2]000), .d(csel[2]0000), .b(vdd), .g(irq));
NEMR4T g256(.s(csel[2]0000), .d(csel[2]00000), .b(vdd), .g(ireset));
NEMR4T g257(.s(csel[2]00000), .d(int_11), .b(vdd), .g(inst[15]));
NEMR4T g258(.s(csel[2]00000), .d(int_16), .b(gnd), .g(inst[15]));
NEMR4T g259(.s(csel[2]00), .d(csel[2]001), .b(gnd), .g(inst[16]));
NEMR4T g260(.s(csel[2]001), .d(csel[2]0010), .b(vdd), .g(irq));
NEMR4T g261(.s(csel[2]0010), .d(csel[2]00100), .b(vdd), .g(ireset));
NEMR4T g262(.s(csel[2]00100), .d(int_13), .b(vdd), .g(inst[15]));
NEMR4T g263(.s(csel[2]00100), .d(int_11), .b(gnd), .g(inst[15]));
NEMR4T g264(.s(csel[2]00), .d(int_16), .b(gnd), .g(ireset));
NEMR4T g265(.s(csel[2]0), .d(csel[2]01), .b(gnd), .g(inst[13]));
NEMR4T g266(.s(csel[2]01), .d(csel[2]011), .b(gnd), .g(inst[16]));
NEMR4T g267(.s(csel[2]011), .d(csel[2]0110), .b(vdd), .g(irq));
NEMR4T g268(.s(csel[2]0110), .d(csel[2]01100), .b(vdd), .g(ireset));
NEMR4T g269(.s(csel[2]01100), .d(int_15), .b(vdd), .g(inst[15]));
NEMR4T g270(.s(csel[2]01), .d(csel[2]0120), .b(vdd), .g(irq));
NEMR4T g271(.s(csel[2]0120), .d(int_34), .b(vdd), .g(ireset));
NEMR4T g272(.s(int_34), .d(int_16), .b(gnd), .g(inst[15]));
NEMR4T g273(.s(csel[2]0120), .d(int_16), .b(vdd), .g(inst[15]));
NEMR4T g274(.s(csel[2]01), .d(int_153), .b(gnd), .g(irq));
NEMR4T g275(.s(int_153), .d(int_35), .b(gnd), .g(ireset));
NEMR4T g276(.s(int_35), .d(int_16), .b(vdd), .g(inst[15]));
NEMR4T g277(.s(csel[2]01), .d(int_34), .b(gnd), .g(ireset));
NEMR4T g278(.s(csel[2]), .d(csel[2]1), .b(gnd), .g(inst[14]));
NEMR4T g279(.s(csel[2]1), .d(csel[2]120), .b(vdd), .g(inst[16]));
NEMR4T g280(.s(csel[2]120), .d(int_35), .b(vdd), .g(irq));
NEMR4T g281(.s(csel[2]120), .d(int_153), .b(gnd), .g(irq));
NEMR4T g282(.s(csel[2]1), .d(csel[2]121), .b(gnd), .g(inst[16]));
NEMR4T g283(.s(csel[2]121), .d(int_154), .b(vdd), .g(irq));
NEMR4T g284(.s(int_154), .d(int_36), .b(vdd), .g(ireset));
NEMR4T g285(.s(int_36), .d(int_13), .b(vdd), .g(inst[15]));
NEMR4T g286(.s(csel[2]121), .d(int_35), .b(gnd), .g(ireset));
NEMR4T g287(.s(csel[2]1), .d(int_37), .b(vdd), .g(irq));
NEMR4T g288(.s(int_37), .d(int_34), .b(vdd), .g(ireset));
NEMR4T g289(.s(csel[2]1), .d(int_34), .b(gnd), .g(ireset));
NEMR4T g290(.s(csel[2]), .d(csel[2]220), .b(vdd), .g(inst[16]));
NEMR4T g291(.s(csel[2]220), .d(csel[2]2200), .b(vdd), .g(irq));
NEMR4T g292(.s(csel[2]2200), .d(int_38), .b(vdd), .g(ireset));
NEMR4T g293(.s(int_38), .d(int_12), .b(vdd), .g(inst[15]));
NEMR4T g294(.s(csel[2]), .d(int_39), .b(vdd), .g(irq));
NEMR4T g295(.s(int_39), .d(int_12), .b(gnd), .g(inst[15]));
NEMR4T g296(.s(csel[2]), .d(int_40), .b(gnd), .g(irq));
NEMR4T g297(.s(int_40), .d(int_13), .b(vdd), .g(ireset));
NEMR4T g298(.s(int_40), .d(int_39), .b(gnd), .g(ireset));
NEMR4T g299(.s(csel[2]), .d(int_38), .b(gnd), .g(ireset));
NEMR4T g300(.s(wsel[0]), .d(wsel[0]0), .b(vdd), .g(inst[15]));
NEMR4T g301(.s(wsel[0]0), .d(int_41), .b(vdd), .g(inst[14]));
NEMR4T g302(.s(int_41), .d(gnd), .b(vdd), .g(inst[17]));
NEMR4T g303(.s(int_41), .d(vdd), .b(gnd), .g(inst[17]));
NEMR4T g304(.s(wsel[0]0), .d(wsel[0]01), .b(gnd), .g(inst[14]));
NEMR4T g305(.s(wsel[0]01), .d(int_0), .b(vdd), .g(inst[13]));
NEMR4T g306(.s(wsel[0]01), .d(int_41), .b(gnd), .g(inst[13]));
NEMR4T g307(.s(wsel[0]), .d(int_41), .b(gnd), .g(inst[15]));
NEMR4T g308(.s(wsel[1]), .d(wsel[1]0), .b(vdd), .g(inst[15]));
NEMR4T g309(.s(wsel[1]0), .d(gnd), .b(vdd), .g(inst[14]));
NEMR4T g310(.s(wsel[1]0), .d(vdd), .b(gnd), .g(inst[14]));
NEMR4T g311(.s(wsel[1]), .d(int_13), .b(gnd), .g(inst[15]));
NEMR4T g312(.s(pcsel[1]), .d(pcsel[1]0), .b(vdd), .g(inst[12]));
NEMR4T g313(.s(pcsel[1]0), .d(pcsel[1]00), .b(vdd), .g(z));
NEMR4T g314(.s(pcsel[1]00), .d(pcsel[1]000), .b(vdd), .g(c));
NEMR4T g315(.s(pcsel[1]000), .d(int_225), .b(vdd), .g(inst[10]));
NEMR4T g316(.s(int_225), .d(int_201), .b(vdd), .g(inst[14]));
NEMR4T g317(.s(int_201), .d(int_156), .b(gnd), .g(inst[13]));
NEMR4T g318(.s(int_156), .d(int_155), .b(vdd), .g(inst[16]));
NEMR4T g319(.s(int_155), .d(int_42), .b(vdd), .g(inst[15]));
NEMR4T g320(.s(int_42), .d(int_1), .b(vdd), .g(irq));
NEMR4T g321(.s(int_42), .d(int_2), .b(gnd), .g(irq));
NEMR4T g322(.s(int_42), .d(vdd), .b(gnd), .g(ireset));
NEMR4T g323(.s(int_155), .d(int_43), .b(gnd), .g(inst[15]));
NEMR4T g324(.s(int_43), .d(int_42), .b(vdd), .g(inst[17]));
NEMR4T g325(.s(int_43), .d(int_0), .b(gnd), .g(inst[17]));
NEMR4T g326(.s(int_156), .d(int_42), .b(gnd), .g(inst[16]));
NEMR4T g327(.s(pcsel[1]00), .d(pcsel[1]001), .b(gnd), .g(c));
NEMR4T g328(.s(pcsel[1]001), .d(int_159), .b(vdd), .g(inst[11]));
NEMR4T g329(.s(int_159), .d(int_158), .b(vdd), .g(inst[14]));
NEMR4T g330(.s(int_158), .d(int_157), .b(vdd), .g(inst[13]));
NEMR4T g331(.s(int_157), .d(int_42), .b(vdd), .g(inst[16]));
NEMR4T g332(.s(int_157), .d(int_155), .b(gnd), .g(inst[16]));
NEMR4T g333(.s(int_158), .d(int_156), .b(gnd), .g(inst[13]));
NEMR4T g334(.s(int_159), .d(int_42), .b(gnd), .g(inst[14]));
NEMR4T g335(.s(pcsel[1]0), .d(pcsel[1]01), .b(gnd), .g(z));
NEMR4T g336(.s(pcsel[1]01), .d(pcsel[1]010), .b(vdd), .g(c));
NEMR4T g337(.s(pcsel[1]010), .d(int_159), .b(gnd), .g(inst[11]));
NEMR4T g338(.s(pcsel[1]01), .d(int_49), .b(vdd), .g(inst[11]));
NEMR4T g339(.s(int_49), .d(int_159), .b(gnd), .g(inst[10]));
NEMR4T g340(.s(pcsel[1]0), .d(pcsel[1]021), .b(gnd), .g(c));
NEMR4T g341(.s(pcsel[1]021), .d(int_49), .b(gnd), .g(inst[11]));
NEMR4T g342(.s(pcsel[1]), .d(pcsel[1]1), .b(gnd), .g(inst[12]));
NEMR4T g343(.s(pcsel[1]1), .d(pcsel[1]10), .b(vdd), .g(z));
NEMR4T g344(.s(pcsel[1]10), .d(pcsel[1]100), .b(vdd), .g(c));
NEMR4T g345(.s(pcsel[1]100), .d(int_160), .b(vdd), .g(inst[10]));
NEMR4T g346(.s(int_160), .d(int_50), .b(vdd), .g(inst[14]));
NEMR4T g347(.s(int_50), .d(int_42), .b(gnd), .g(inst[13]));
NEMR4T g348(.s(pcsel[1]10), .d(pcsel[1]101), .b(gnd), .g(c));
NEMR4T g349(.s(pcsel[1]101), .d(int_202), .b(vdd), .g(inst[11]));
NEMR4T g350(.s(int_202), .d(int_52), .b(vdd), .g(inst[10]));
NEMR4T g351(.s(int_52), .d(int_51), .b(vdd), .g(inst[14]));
NEMR4T g352(.s(int_51), .d(int_157), .b(vdd), .g(inst[13]));
NEMR4T g353(.s(int_51), .d(int_42), .b(gnd), .g(inst[13]));
NEMR4T g354(.s(int_52), .d(int_42), .b(gnd), .g(inst[14]));
NEMR4T g355(.s(int_202), .d(int_225), .b(gnd), .g(inst[10]));
NEMR4T g356(.s(pcsel[1]1), .d(pcsel[1]11), .b(gnd), .g(z));
NEMR4T g357(.s(pcsel[1]11), .d(pcsel[1]110), .b(vdd), .g(c));
NEMR4T g358(.s(pcsel[1]110), .d(int_202), .b(gnd), .g(inst[11]));
NEMR4T g359(.s(pcsel[1]110), .d(int_56), .b(gnd), .g(inst[10]));
NEMR4T g360(.s(int_56), .d(int_55), .b(vdd), .g(inst[14]));
NEMR4T g361(.s(int_55), .d(int_157), .b(vdd), .g(inst[13]));
NEMR4T g362(.s(int_56), .d(int_42), .b(gnd), .g(inst[14]));
NEMR4T g363(.s(pcsel[1]11), .d(int_162), .b(vdd), .g(inst[11]));
NEMR4T g364(.s(int_162), .d(int_160), .b(gnd), .g(inst[10]));
NEMR4T g365(.s(pcsel[1]1), .d(pcsel[1]121), .b(gnd), .g(c));
NEMR4T g366(.s(pcsel[1]121), .d(int_162), .b(gnd), .g(inst[11]));
NEMR4T g367(.s(pcsel[1]121), .d(int_56), .b(gnd), .g(inst[10]));
NEMR4T g368(.s(pcsel[1]), .d(pcsel[1]20), .b(vdd), .g(z));
NEMR4T g369(.s(pcsel[1]20), .d(pcsel[1]200), .b(vdd), .g(c));
NEMR4T g370(.s(pcsel[1]200), .d(int_225), .b(gnd), .g(inst[10]));
NEMR4T g371(.s(pcsel[1]200), .d(int_55), .b(vdd), .g(inst[14]));
NEMR4T g372(.s(pcsel[1]200), .d(int_42), .b(gnd), .g(inst[14]));
NEMR4T g373(.s(pcsel[1]), .d(pcsel[1]21), .b(gnd), .g(z));
NEMR4T g374(.s(pcsel[1]21), .d(int_58), .b(vdd), .g(inst[11]));
NEMR4T g375(.s(int_58), .d(int_159), .b(vdd), .g(inst[10]));
NEMR4T g376(.s(pcsel[1]), .d(pcsel[1]221), .b(gnd), .g(c));
NEMR4T g377(.s(pcsel[1]221), .d(int_58), .b(gnd), .g(inst[11]));
NEMR4T g378(.s(pcsel[0]), .d(pcsel[0]0), .b(vdd), .g(inst[12]));
NEMR4T g379(.s(pcsel[0]0), .d(pcsel[0]00), .b(vdd), .g(z));
NEMR4T g380(.s(pcsel[0]00), .d(pcsel[0]000), .b(vdd), .g(c));
NEMR4T g381(.s(pcsel[0]000), .d(int_163), .b(vdd), .g(inst[10]));
NEMR4T g382(.s(int_163), .d(int_61), .b(gnd), .g(inst[17]));
NEMR4T g383(.s(int_61), .d(int_60), .b(vdd), .g(inst[15]));
NEMR4T g384(.s(int_60), .d(int_59), .b(vdd), .g(inst[13]));
NEMR4T g385(.s(int_59), .d(int_42), .b(vdd), .g(inst[16]));
NEMR4T g386(.s(int_59), .d(int_0), .b(gnd), .g(inst[16]));
NEMR4T g387(.s(int_60), .d(int_42), .b(gnd), .g(inst[13]));
NEMR4T g388(.s(int_61), .d(int_42), .b(gnd), .g(inst[15]));
NEMR4T g389(.s(pcsel[0]00), .d(pcsel[0]001), .b(gnd), .g(c));
NEMR4T g390(.s(pcsel[0]001), .d(int_62), .b(vdd), .g(inst[11]));
NEMR4T g391(.s(int_62), .d(int_42), .b(vdd), .g(inst[17]));
NEMR4T g392(.s(int_62), .d(int_61), .b(gnd), .g(inst[17]));
NEMR4T g393(.s(pcsel[0]0), .d(pcsel[0]01), .b(gnd), .g(z));
NEMR4T g394(.s(pcsel[0]01), .d(pcsel[0]010), .b(vdd), .g(c));
NEMR4T g395(.s(pcsel[0]010), .d(int_62), .b(gnd), .g(inst[11]));
NEMR4T g396(.s(pcsel[0]01), .d(int_63), .b(vdd), .g(inst[11]));
NEMR4T g397(.s(int_63), .d(int_62), .b(gnd), .g(inst[10]));
NEMR4T g398(.s(pcsel[0]0), .d(pcsel[0]021), .b(gnd), .g(c));
NEMR4T g399(.s(pcsel[0]021), .d(int_63), .b(gnd), .g(inst[11]));
NEMR4T g400(.s(pcsel[0]), .d(pcsel[0]1), .b(gnd), .g(inst[12]));
NEMR4T g401(.s(pcsel[0]1), .d(pcsel[0]10), .b(vdd), .g(z));
NEMR4T g402(.s(pcsel[0]10), .d(pcsel[0]100), .b(vdd), .g(c));
NEMR4T g403(.s(pcsel[0]100), .d(int_64), .b(vdd), .g(inst[10]));
NEMR4T g404(.s(int_64), .d(int_42), .b(gnd), .g(inst[17]));
NEMR4T g405(.s(pcsel[0]10), .d(pcsel[0]101), .b(gnd), .g(c));
NEMR4T g406(.s(pcsel[0]101), .d(int_164), .b(vdd), .g(inst[11]));
NEMR4T g407(.s(int_164), .d(int_42), .b(vdd), .g(inst[10]));
NEMR4T g408(.s(int_164), .d(int_163), .b(gnd), .g(inst[10]));
NEMR4T g409(.s(pcsel[0]1), .d(pcsel[0]11), .b(gnd), .g(z));
NEMR4T g410(.s(pcsel[0]11), .d(pcsel[0]110), .b(vdd), .g(c));
NEMR4T g411(.s(pcsel[0]110), .d(int_164), .b(gnd), .g(inst[11]));
NEMR4T g412(.s(pcsel[0]110), .d(int_66), .b(gnd), .g(inst[10]));
NEMR4T g413(.s(int_66), .d(int_42), .b(vdd), .g(inst[17]));
NEMR4T g414(.s(pcsel[0]11), .d(int_67), .b(vdd), .g(inst[11]));
NEMR4T g415(.s(int_67), .d(int_64), .b(gnd), .g(inst[10]));
NEMR4T g416(.s(pcsel[0]1), .d(pcsel[0]121), .b(gnd), .g(c));
NEMR4T g417(.s(pcsel[0]121), .d(int_67), .b(gnd), .g(inst[11]));
NEMR4T g418(.s(pcsel[0]121), .d(int_66), .b(gnd), .g(inst[10]));
NEMR4T g419(.s(pcsel[0]), .d(pcsel[0]20), .b(vdd), .g(z));
NEMR4T g420(.s(pcsel[0]20), .d(pcsel[0]200), .b(vdd), .g(c));
NEMR4T g421(.s(pcsel[0]200), .d(int_163), .b(gnd), .g(inst[10]));
NEMR4T g422(.s(pcsel[0]200), .d(int_42), .b(vdd), .g(inst[17]));
NEMR4T g423(.s(pcsel[0]), .d(pcsel[0]21), .b(gnd), .g(z));
NEMR4T g424(.s(pcsel[0]21), .d(int_68), .b(vdd), .g(inst[11]));
NEMR4T g425(.s(int_68), .d(int_62), .b(vdd), .g(inst[10]));
NEMR4T g426(.s(pcsel[0]), .d(pcsel[0]221), .b(gnd), .g(c));
NEMR4T g427(.s(pcsel[0]221), .d(int_68), .b(gnd), .g(inst[11]));
NEMR4T g428(.s(stsel[0]), .d(stsel[0]0), .b(vdd), .g(inst[12]));
NEMR4T g429(.s(stsel[0]0), .d(stsel[0]00), .b(vdd), .g(z));
NEMR4T g430(.s(stsel[0]00), .d(stsel[0]000), .b(vdd), .g(c));
NEMR4T g431(.s(stsel[0]000), .d(int_206), .b(vdd), .g(inst[10]));
NEMR4T g432(.s(int_206), .d(int_205), .b(gnd), .g(inst[17]));
NEMR4T g433(.s(int_205), .d(int_204), .b(vdd), .g(inst[15]));
NEMR4T g434(.s(int_204), .d(int_203), .b(vdd), .g(inst[14]));
NEMR4T g435(.s(int_203), .d(int_165), .b(vdd), .g(inst[13]));
NEMR4T g436(.s(int_165), .d(int_69), .b(gnd), .g(inst[16]));
NEMR4T g437(.s(int_69), .d(vdd), .b(vdd), .g(ireset));
NEMR4T g438(.s(int_69), .d(gnd), .b(gnd), .g(ireset));
NEMR4T g439(.s(int_204), .d(int_70), .b(gnd), .g(inst[14]));
NEMR4T g440(.s(int_70), .d(int_1), .b(vdd), .g(irq));
NEMR4T g441(.s(int_70), .d(int_2), .b(gnd), .g(irq));
NEMR4T g442(.s(int_70), .d(gnd), .b(gnd), .g(ireset));
NEMR4T g443(.s(int_205), .d(int_167), .b(gnd), .g(inst[15]));
NEMR4T g444(.s(int_167), .d(int_166), .b(vdd), .g(inst[14]));
NEMR4T g445(.s(int_166), .d(int_71), .b(vdd), .g(inst[13]));
NEMR4T g446(.s(int_71), .d(int_70), .b(vdd), .g(inst[16]));
NEMR4T g447(.s(int_167), .d(int_73), .b(gnd), .g(inst[14]));
NEMR4T g448(.s(int_73), .d(int_72), .b(gnd), .g(inst[13]));
NEMR4T g449(.s(int_72), .d(int_70), .b(gnd), .g(inst[16]));
NEMR4T g450(.s(int_73), .d(int_70), .b(vdd), .g(inst[16]));
NEMR4T g451(.s(int_167), .d(int_72), .b(vdd), .g(inst[13]));
NEMR4T g452(.s(int_206), .d(int_168), .b(vdd), .g(inst[15]));
NEMR4T g453(.s(int_168), .d(int_166), .b(vdd), .g(inst[14]));
NEMR4T g454(.s(stsel[0]00), .d(stsel[0]001), .b(gnd), .g(c));
NEMR4T g455(.s(stsel[0]001), .d(int_172), .b(vdd), .g(inst[11]));
NEMR4T g456(.s(int_172), .d(int_75), .b(vdd), .g(inst[17]));
NEMR4T g457(.s(int_75), .d(int_73), .b(gnd), .g(inst[14]));
NEMR4T g458(.s(int_75), .d(int_72), .b(vdd), .g(inst[13]));
NEMR4T g459(.s(int_172), .d(int_171), .b(gnd), .g(inst[17]));
NEMR4T g460(.s(int_171), .d(int_204), .b(vdd), .g(inst[15]));
NEMR4T g461(.s(int_171), .d(int_75), .b(gnd), .g(inst[15]));
NEMR4T g462(.s(int_172), .d(int_168), .b(gnd), .g(inst[15]));
NEMR4T g463(.s(int_172), .d(int_78), .b(vdd), .g(inst[14]));
NEMR4T g464(.s(int_78), .d(int_70), .b(gnd), .g(inst[13]));
NEMR4T g465(.s(stsel[0]0), .d(stsel[0]01), .b(gnd), .g(z));
NEMR4T g466(.s(stsel[0]01), .d(stsel[0]010), .b(vdd), .g(c));
NEMR4T g467(.s(stsel[0]010), .d(int_172), .b(gnd), .g(inst[11]));
NEMR4T g468(.s(stsel[0]01), .d(int_207), .b(vdd), .g(inst[11]));
NEMR4T g469(.s(int_207), .d(int_173), .b(gnd), .g(inst[10]));
NEMR4T g470(.s(int_173), .d(int_75), .b(vdd), .g(inst[17]));
NEMR4T g471(.s(int_173), .d(int_171), .b(gnd), .g(inst[17]));
NEMR4T g472(.s(int_173), .d(int_82), .b(vdd), .g(inst[14]));
NEMR4T g473(.s(int_82), .d(int_71), .b(vdd), .g(inst[13]));
NEMR4T g474(.s(int_82), .d(int_70), .b(gnd), .g(inst[13]));
NEMR4T g475(.s(stsel[0]0), .d(stsel[0]021), .b(gnd), .g(c));
NEMR4T g476(.s(stsel[0]021), .d(int_207), .b(gnd), .g(inst[11]));
NEMR4T g477(.s(stsel[0]), .d(stsel[0]1), .b(gnd), .g(inst[12]));
NEMR4T g478(.s(stsel[0]1), .d(stsel[0]10), .b(vdd), .g(z));
NEMR4T g479(.s(stsel[0]10), .d(stsel[0]100), .b(vdd), .g(c));
NEMR4T g480(.s(stsel[0]100), .d(stsel[0]10020), .b(vdd), .g(inst[10]));
NEMR4T g481(.s(stsel[0]10020), .d(int_84), .b(vdd), .g(inst[17]));
NEMR4T g482(.s(int_84), .d(int_168), .b(vdd), .g(inst[15]));
NEMR4T g483(.s(stsel[0]10020), .d(int_167), .b(gnd), .g(inst[17]));
NEMR4T g484(.s(stsel[0]10), .d(stsel[0]101), .b(gnd), .g(c));
NEMR4T g485(.s(stsel[0]101), .d(int_208), .b(vdd), .g(inst[11]));
NEMR4T g486(.s(int_208), .d(int_86), .b(vdd), .g(inst[10]));
NEMR4T g487(.s(int_86), .d(int_168), .b(gnd), .g(inst[15]));
NEMR4T g488(.s(int_86), .d(int_78), .b(vdd), .g(inst[14]));
NEMR4T g489(.s(int_86), .d(int_73), .b(gnd), .g(inst[14]));
NEMR4T g490(.s(int_86), .d(int_72), .b(vdd), .g(inst[13]));
NEMR4T g491(.s(int_208), .d(int_174), .b(gnd), .g(inst[10]));
NEMR4T g492(.s(int_174), .d(int_87), .b(gnd), .g(inst[17]));
NEMR4T g493(.s(int_87), .d(int_204), .b(vdd), .g(inst[15]));
NEMR4T g494(.s(int_87), .d(int_167), .b(gnd), .g(inst[15]));
NEMR4T g495(.s(int_87), .d(int_78), .b(vdd), .g(inst[14]));
NEMR4T g496(.s(stsel[0]1), .d(stsel[0]11), .b(gnd), .g(z));
NEMR4T g497(.s(stsel[0]11), .d(stsel[0]110), .b(vdd), .g(c));
NEMR4T g498(.s(stsel[0]110), .d(int_208), .b(gnd), .g(inst[11]));
NEMR4T g499(.s(stsel[0]110), .d(int_88), .b(gnd), .g(inst[10]));
NEMR4T g500(.s(int_88), .d(int_86), .b(vdd), .g(inst[17]));
NEMR4T g501(.s(stsel[0]11), .d(int_209), .b(vdd), .g(inst[11]));
NEMR4T g502(.s(int_209), .d(int_175), .b(gnd), .g(inst[10]));
NEMR4T g503(.s(int_175), .d(int_84), .b(vdd), .g(inst[17]));
NEMR4T g504(.s(int_175), .d(int_89), .b(gnd), .g(inst[17]));
NEMR4T g505(.s(int_89), .d(int_82), .b(vdd), .g(inst[14]));
NEMR4T g506(.s(int_89), .d(int_73), .b(gnd), .g(inst[14]));
NEMR4T g507(.s(int_89), .d(int_72), .b(vdd), .g(inst[13]));
NEMR4T g508(.s(stsel[0]1), .d(stsel[0]121), .b(gnd), .g(c));
NEMR4T g509(.s(stsel[0]121), .d(int_209), .b(gnd), .g(inst[11]));
NEMR4T g510(.s(stsel[0]121), .d(int_88), .b(gnd), .g(inst[10]));
NEMR4T g511(.s(stsel[0]), .d(stsel[0]20), .b(vdd), .g(z));
NEMR4T g512(.s(stsel[0]20), .d(stsel[0]200), .b(vdd), .g(c));
NEMR4T g513(.s(stsel[0]200), .d(int_206), .b(gnd), .g(inst[10]));
NEMR4T g514(.s(stsel[0]200), .d(stsel[0]200220), .b(vdd), .g(inst[17]));
NEMR4T g515(.s(stsel[0]200220), .d(int_168), .b(gnd), .g(inst[15]));
NEMR4T g516(.s(stsel[0]200220), .d(int_73), .b(gnd), .g(inst[14]));
NEMR4T g517(.s(stsel[0]200220), .d(int_72), .b(vdd), .g(inst[13]));
NEMR4T g518(.s(stsel[0]200), .d(int_78), .b(vdd), .g(inst[14]));
NEMR4T g519(.s(stsel[0]20), .d(stsel[0]201), .b(gnd), .g(c));
NEMR4T g520(.s(stsel[0]201), .d(int_84), .b(vdd), .g(inst[11]));
NEMR4T g521(.s(stsel[0]), .d(stsel[0]21), .b(gnd), .g(z));
NEMR4T g522(.s(stsel[0]21), .d(stsel[0]210), .b(vdd), .g(c));
NEMR4T g523(.s(stsel[0]210), .d(int_84), .b(gnd), .g(inst[11]));
NEMR4T g524(.s(stsel[0]21), .d(int_90), .b(vdd), .g(inst[11]));
NEMR4T g525(.s(int_90), .d(int_173), .b(vdd), .g(inst[10]));
NEMR4T g526(.s(stsel[0]), .d(stsel[0]221), .b(gnd), .g(c));
NEMR4T g527(.s(stsel[0]221), .d(int_90), .b(gnd), .g(inst[11]));
NEMR4T g528(.s(stsel[1]), .d(stsel[1]0), .b(vdd), .g(inst[12]));
NEMR4T g529(.s(stsel[1]0), .d(stsel[1]00), .b(vdd), .g(z));
NEMR4T g530(.s(stsel[1]00), .d(stsel[1]000), .b(vdd), .g(c));
NEMR4T g531(.s(stsel[1]000), .d(int_210), .b(vdd), .g(inst[10]));
NEMR4T g532(.s(int_210), .d(int_179), .b(vdd), .g(inst[14]));
NEMR4T g533(.s(int_179), .d(int_178), .b(gnd), .g(inst[13]));
NEMR4T g534(.s(int_178), .d(int_177), .b(vdd), .g(inst[16]));
NEMR4T g535(.s(int_177), .d(int_176), .b(vdd), .g(irq));
NEMR4T g536(.s(int_176), .d(int_91), .b(vdd), .g(ireset));
NEMR4T g537(.s(int_91), .d(int_11), .b(gnd), .g(inst[15]));
NEMR4T g538(.s(int_177), .d(int_92), .b(gnd), .g(irq));
NEMR4T g539(.s(int_92), .d(int_39), .b(gnd), .g(ireset));
NEMR4T g540(.s(int_178), .d(int_93), .b(gnd), .g(inst[16]));
NEMR4T g541(.s(int_93), .d(int_37), .b(vdd), .g(irq));
NEMR4T g542(.s(int_179), .d(int_94), .b(gnd), .g(inst[16]));
NEMR4T g543(.s(int_94), .d(int_92), .b(gnd), .g(irq));
NEMR4T g544(.s(stsel[1]00), .d(stsel[1]001), .b(gnd), .g(c));
NEMR4T g545(.s(stsel[1]001), .d(int_213), .b(vdd), .g(inst[11]));
NEMR4T g546(.s(int_213), .d(int_212), .b(vdd), .g(inst[14]));
NEMR4T g547(.s(int_212), .d(int_211), .b(vdd), .g(inst[13]));
NEMR4T g548(.s(int_211), .d(int_93), .b(vdd), .g(inst[16]));
NEMR4T g549(.s(int_211), .d(int_180), .b(gnd), .g(inst[16]));
NEMR4T g550(.s(int_180), .d(int_176), .b(vdd), .g(irq));
NEMR4T g551(.s(int_212), .d(int_97), .b(gnd), .g(inst[13]));
NEMR4T g552(.s(int_97), .d(int_180), .b(vdd), .g(inst[16]));
NEMR4T g553(.s(int_97), .d(int_93), .b(gnd), .g(inst[16]));
NEMR4T g554(.s(int_213), .d(int_93), .b(gnd), .g(inst[14]));
NEMR4T g555(.s(int_213), .d(int_98), .b(vdd), .g(irq));
NEMR4T g556(.s(int_98), .d(int_36), .b(vdd), .g(ireset));
NEMR4T g557(.s(int_98), .d(int_12), .b(gnd), .g(inst[15]));
NEMR4T g558(.s(int_213), .d(int_40), .b(gnd), .g(irq));
NEMR4T g559(.s(int_213), .d(int_99), .b(gnd), .g(ireset));
NEMR4T g560(.s(int_99), .d(int_12), .b(vdd), .g(inst[15]));
NEMR4T g561(.s(int_99), .d(gnd), .b(gnd), .g(inst[17]));
NEMR4T g562(.s(stsel[1]0), .d(stsel[1]01), .b(gnd), .g(z));
NEMR4T g563(.s(stsel[1]01), .d(stsel[1]010), .b(vdd), .g(c));
NEMR4T g564(.s(stsel[1]010), .d(int_213), .b(gnd), .g(inst[11]));
NEMR4T g565(.s(stsel[1]01), .d(int_214), .b(vdd), .g(inst[11]));
NEMR4T g566(.s(int_214), .d(int_181), .b(gnd), .g(inst[10]));
NEMR4T g567(.s(int_181), .d(int_102), .b(vdd), .g(inst[14]));
NEMR4T g568(.s(int_102), .d(int_101), .b(vdd), .g(inst[13]));
NEMR4T g569(.s(int_101), .d(int_93), .b(vdd), .g(inst[16]));
NEMR4T g570(.s(int_101), .d(int_180), .b(gnd), .g(inst[16]));
NEMR4T g571(.s(int_101), .d(int_98), .b(vdd), .g(irq));
NEMR4T g572(.s(int_101), .d(int_40), .b(gnd), .g(irq));
NEMR4T g573(.s(int_101), .d(int_99), .b(gnd), .g(ireset));
NEMR4T g574(.s(int_102), .d(int_97), .b(gnd), .g(inst[13]));
NEMR4T g575(.s(int_181), .d(int_105), .b(gnd), .g(inst[14]));
NEMR4T g576(.s(int_105), .d(int_104), .b(vdd), .g(irq));
NEMR4T g577(.s(int_104), .d(int_103), .b(vdd), .g(ireset));
NEMR4T g578(.s(int_103), .d(int_13), .b(vdd), .g(inst[15]));
NEMR4T g579(.s(int_103), .d(int_16), .b(gnd), .g(inst[15]));
NEMR4T g580(.s(int_104), .d(int_12), .b(gnd), .g(inst[15]));
NEMR4T g581(.s(int_105), .d(int_40), .b(gnd), .g(irq));
NEMR4T g582(.s(int_105), .d(int_99), .b(gnd), .g(ireset));
NEMR4T g583(.s(stsel[1]0), .d(stsel[1]021), .b(gnd), .g(c));
NEMR4T g584(.s(stsel[1]021), .d(int_214), .b(gnd), .g(inst[11]));
NEMR4T g585(.s(stsel[1]), .d(stsel[1]1), .b(gnd), .g(inst[12]));
NEMR4T g586(.s(stsel[1]1), .d(stsel[1]10), .b(vdd), .g(z));
NEMR4T g587(.s(stsel[1]10), .d(stsel[1]100), .b(vdd), .g(c));
NEMR4T g588(.s(stsel[1]100), .d(stsel[1]10020), .b(vdd), .g(inst[10]));
NEMR4T g589(.s(stsel[1]10020), .d(stsel[1]100200), .b(vdd), .g(inst[14]));
NEMR4T g590(.s(stsel[1]100200), .d(int_107), .b(vdd), .g(inst[13]));
NEMR4T g591(.s(int_107), .d(int_94), .b(gnd), .g(inst[16]));
NEMR4T g592(.s(stsel[1]100200), .d(int_108), .b(gnd), .g(inst[13]));
NEMR4T g593(.s(int_108), .d(int_37), .b(vdd), .g(irq));
NEMR4T g594(.s(int_108), .d(int_92), .b(gnd), .g(irq));
NEMR4T g595(.s(stsel[1]10), .d(stsel[1]101), .b(gnd), .g(c));
NEMR4T g596(.s(stsel[1]101), .d(int_215), .b(vdd), .g(inst[11]));
NEMR4T g597(.s(int_215), .d(int_110), .b(vdd), .g(inst[10]));
NEMR4T g598(.s(int_110), .d(int_109), .b(vdd), .g(inst[14]));
NEMR4T g599(.s(int_109), .d(int_211), .b(vdd), .g(inst[13]));
NEMR4T g600(.s(int_109), .d(int_93), .b(gnd), .g(inst[13]));
NEMR4T g601(.s(int_110), .d(int_93), .b(gnd), .g(inst[14]));
NEMR4T g602(.s(int_110), .d(int_98), .b(vdd), .g(irq));
NEMR4T g603(.s(int_110), .d(int_40), .b(gnd), .g(irq));
NEMR4T g604(.s(int_110), .d(int_99), .b(gnd), .g(ireset));
NEMR4T g605(.s(int_215), .d(int_182), .b(gnd), .g(inst[10]));
NEMR4T g606(.s(int_182), .d(int_113), .b(vdd), .g(inst[14]));
NEMR4T g607(.s(int_113), .d(int_112), .b(gnd), .g(inst[13]));
NEMR4T g608(.s(int_112), .d(int_177), .b(vdd), .g(inst[16]));
NEMR4T g609(.s(int_112), .d(int_93), .b(gnd), .g(inst[16]));
NEMR4T g610(.s(int_112), .d(int_98), .b(vdd), .g(irq));
NEMR4T g611(.s(int_112), .d(int_145), .b(gnd), .g(irq));
NEMR4T g612(.s(int_112), .d(int_99), .b(gnd), .g(ireset));
NEMR4T g613(.s(int_113), .d(int_94), .b(gnd), .g(inst[16]));
NEMR4T g614(.s(stsel[1]1), .d(stsel[1]11), .b(gnd), .g(z));
NEMR4T g615(.s(stsel[1]11), .d(stsel[1]110), .b(vdd), .g(c));
NEMR4T g616(.s(stsel[1]110), .d(int_215), .b(gnd), .g(inst[11]));
NEMR4T g617(.s(stsel[1]110), .d(int_184), .b(gnd), .g(inst[10]));
NEMR4T g618(.s(int_184), .d(int_183), .b(vdd), .g(inst[14]));
NEMR4T g619(.s(int_183), .d(int_114), .b(vdd), .g(inst[13]));
NEMR4T g620(.s(int_114), .d(int_108), .b(vdd), .g(inst[16]));
NEMR4T g621(.s(int_114), .d(int_180), .b(gnd), .g(inst[16]));
NEMR4T g622(.s(int_114), .d(int_98), .b(vdd), .g(irq));
NEMR4T g623(.s(int_114), .d(int_145), .b(gnd), .g(irq));
NEMR4T g624(.s(int_114), .d(int_99), .b(gnd), .g(ireset));
NEMR4T g625(.s(int_184), .d(int_105), .b(gnd), .g(inst[14]));
NEMR4T g626(.s(stsel[1]11), .d(int_216), .b(vdd), .g(inst[11]));
NEMR4T g627(.s(int_216), .d(int_185), .b(gnd), .g(inst[10]));
NEMR4T g628(.s(int_185), .d(int_115), .b(vdd), .g(inst[14]));
NEMR4T g629(.s(int_115), .d(int_107), .b(vdd), .g(inst[13]));
NEMR4T g630(.s(int_115), .d(int_93), .b(gnd), .g(inst[13]));
NEMR4T g631(.s(stsel[1]1), .d(stsel[1]121), .b(gnd), .g(c));
NEMR4T g632(.s(stsel[1]121), .d(int_216), .b(gnd), .g(inst[11]));
NEMR4T g633(.s(stsel[1]121), .d(int_184), .b(gnd), .g(inst[10]));
NEMR4T g634(.s(stsel[1]), .d(stsel[1]20), .b(vdd), .g(z));
NEMR4T g635(.s(stsel[1]20), .d(stsel[1]200), .b(vdd), .g(c));
NEMR4T g636(.s(stsel[1]200), .d(int_210), .b(gnd), .g(inst[10]));
NEMR4T g637(.s(stsel[1]200), .d(stsel[1]200220), .b(vdd), .g(inst[14]));
NEMR4T g638(.s(stsel[1]200220), .d(stsel[1]2002200), .b(vdd), .g(inst[13]));
NEMR4T g639(.s(stsel[1]2002200), .d(int_108), .b(vdd), .g(inst[16]));
NEMR4T g640(.s(stsel[1]2002200), .d(int_180), .b(gnd), .g(inst[16]));
NEMR4T g641(.s(stsel[1]200), .d(int_108), .b(gnd), .g(inst[14]));
NEMR4T g642(.s(stsel[1]200), .d(int_98), .b(vdd), .g(irq));
NEMR4T g643(.s(stsel[1]200), .d(int_145), .b(gnd), .g(irq));
NEMR4T g644(.s(stsel[1]200), .d(int_99), .b(gnd), .g(ireset));
NEMR4T g645(.s(stsel[1]), .d(stsel[1]21), .b(gnd), .g(z));
NEMR4T g646(.s(stsel[1]21), .d(int_217), .b(vdd), .g(inst[11]));
NEMR4T g647(.s(int_217), .d(int_181), .b(vdd), .g(inst[10]));
NEMR4T g648(.s(int_217), .d(int_186), .b(vdd), .g(inst[14]));
NEMR4T g649(.s(int_186), .d(int_116), .b(gnd), .g(inst[13]));
NEMR4T g650(.s(int_116), .d(int_98), .b(vdd), .g(irq));
NEMR4T g651(.s(int_116), .d(int_40), .b(gnd), .g(irq));
NEMR4T g652(.s(int_116), .d(int_99), .b(gnd), .g(ireset));
NEMR4T g653(.s(stsel[1]), .d(stsel[1]221), .b(gnd), .g(c));
NEMR4T g654(.s(stsel[1]221), .d(int_217), .b(gnd), .g(inst[11]));
NEMR4T g655(.s(read_strobe), .d(read_strobe0), .b(vdd), .g(irq));
NEMR4T g656(.s(read_strobe0), .d(read_strobe00), .b(vdd), .g(ireset));
NEMR4T g657(.s(read_strobe00), .d(read_strobe000), .b(vdd), .g(inst[17]));
NEMR4T g658(.s(read_strobe000), .d(read_strobe0000), .b(vdd), .g(inst[13]));
NEMR4T g659(.s(read_strobe0000), .d(read_strobe00000), .b(vdd), .g(inst[16]));
NEMR4T g660(.s(read_strobe00000), .d(int_117), .b(vdd), .g(inst[15]));
NEMR4T g661(.s(int_117), .d(vdd), .b(gnd), .g(inst[14]));
NEMR4T g662(.s(read_strobe00000), .d(int_13), .b(gnd), .g(inst[15]));
NEMR4T g663(.s(read_strobe0000), .d(int_13), .b(gnd), .g(inst[16]));
NEMR4T g664(.s(read_strobe000), .d(int_13), .b(gnd), .g(inst[13]));
NEMR4T g665(.s(read_strobe0), .d(read_strobe01), .b(gnd), .g(ireset));
NEMR4T g666(.s(read_strobe01), .d(int_226), .b(gnd), .g(inst[17]));
NEMR4T g667(.s(int_226), .d(int_218), .b(vdd), .g(inst[13]));
NEMR4T g668(.s(int_218), .d(int_187), .b(vdd), .g(inst[16]));
NEMR4T g669(.s(int_187), .d(int_118), .b(vdd), .g(inst[15]));
NEMR4T g670(.s(int_118), .d(gnd), .b(vdd), .g(inst[14]));
NEMR4T g671(.s(read_strobe0), .d(int_189), .b(gnd), .g(inst[17]));
NEMR4T g672(.s(int_189), .d(int_188), .b(vdd), .g(inst[13]));
NEMR4T g673(.s(int_188), .d(int_187), .b(gnd), .g(inst[16]));
NEMR4T g674(.s(int_189), .d(int_187), .b(gnd), .g(inst[13]));
NEMR4T g675(.s(int_189), .d(int_118), .b(gnd), .g(inst[15]));
NEMR4T g676(.s(int_189), .d(gnd), .b(gnd), .g(inst[14]));
NEMR4T g677(.s(read_strobe), .d(read_strobe1), .b(gnd), .g(irq));
NEMR4T g678(.s(read_strobe1), .d(int_189), .b(vdd), .g(ireset));
NEMR4T g679(.s(read_strobe1), .d(int_120), .b(gnd), .g(ireset));
NEMR4T g680(.s(int_120), .d(int_13), .b(gnd), .g(inst[17]));
NEMR4T g681(.s(read_strobe), .d(int_226), .b(vdd), .g(ireset));
NEMR4T g682(.s(read_strobe), .d(int_121), .b(gnd), .g(ireset));
NEMR4T g683(.s(int_121), .d(int_13), .b(vdd), .g(inst[17]));
NEMR4T g684(.s(write_strobe), .d(write_strobe0), .b(vdd), .g(inst[13]));
NEMR4T g685(.s(write_strobe0), .d(write_strobe00), .b(vdd), .g(inst[16]));
NEMR4T g686(.s(write_strobe00), .d(write_strobe000), .b(vdd), .g(clk));
NEMR4T g687(.s(write_strobe000), .d(write_strobe0000), .b(vdd), .g(irq));
NEMR4T g688(.s(write_strobe0000), .d(write_strobe00000), .b(vdd), .g(ireset));
NEMR4T g689(.s(write_strobe00000), .d(int_13), .b(vdd), .g(inst[15]));
NEMR4T g690(.s(write_strobe00000), .d(write_strobe000001), .b(gnd), .g(inst[15]));
NEMR4T g691(.s(write_strobe000001), .d(int_117), .b(gnd), .g(inst[17]));
NEMR4T g692(.s(write_strobe0000), .d(int_121), .b(gnd), .g(inst[15]));
NEMR4T g693(.s(write_strobe000), .d(int_190), .b(gnd), .g(irq));
NEMR4T g694(.s(int_190), .d(int_13), .b(vdd), .g(ireset));
NEMR4T g695(.s(int_190), .d(int_122), .b(gnd), .g(ireset));
NEMR4T g696(.s(int_122), .d(int_121), .b(gnd), .g(inst[15]));
NEMR4T g697(.s(write_strobe000), .d(int_123), .b(gnd), .g(ireset));
NEMR4T g698(.s(int_123), .d(int_121), .b(vdd), .g(inst[15]));
NEMR4T g699(.s(int_123), .d(int_13), .b(gnd), .g(inst[17]));
NEMR4T g700(.s(write_strobe0), .d(int_221), .b(gnd), .g(inst[16]));
NEMR4T g701(.s(int_221), .d(int_220), .b(vdd), .g(irq));
NEMR4T g702(.s(int_220), .d(int_219), .b(vdd), .g(ireset));
NEMR4T g703(.s(int_219), .d(int_13), .b(vdd), .g(inst[15]));
NEMR4T g704(.s(int_219), .d(int_191), .b(gnd), .g(inst[15]));
NEMR4T g705(.s(int_191), .d(int_124), .b(gnd), .g(inst[17]));
NEMR4T g706(.s(int_124), .d(gnd), .b(gnd), .g(inst[14]));
NEMR4T g707(.s(int_220), .d(int_121), .b(gnd), .g(inst[15]));
NEMR4T g708(.s(int_221), .d(int_190), .b(gnd), .g(irq));
NEMR4T g709(.s(int_221), .d(int_123), .b(gnd), .g(ireset));
NEMR4T g710(.s(write_strobe0), .d(int_222), .b(vdd), .g(irq));
NEMR4T g711(.s(int_222), .d(int_192), .b(vdd), .g(ireset));
NEMR4T g712(.s(int_192), .d(int_126), .b(gnd), .g(inst[15]));
NEMR4T g713(.s(int_126), .d(int_118), .b(gnd), .g(inst[17]));
NEMR4T g714(.s(write_strobe), .d(write_strobe1), .b(gnd), .g(inst[13]));
NEMR4T g715(.s(write_strobe1), .d(write_strobe10), .b(vdd), .g(inst[16]));
NEMR4T g716(.s(write_strobe10), .d(write_strobe101), .b(gnd), .g(clk));
NEMR4T g717(.s(write_strobe101), .d(int_222), .b(vdd), .g(irq));
NEMR4T g718(.s(write_strobe1), .d(write_strobe11), .b(gnd), .g(inst[16]));
NEMR4T g719(.s(write_strobe11), .d(int_129), .b(gnd), .g(clk));
NEMR4T g720(.s(int_129), .d(int_128), .b(vdd), .g(irq));
NEMR4T g721(.s(int_128), .d(int_127), .b(vdd), .g(ireset));
NEMR4T g722(.s(int_127), .d(int_13), .b(vdd), .g(inst[15]));
NEMR4T g723(.s(int_127), .d(int_120), .b(gnd), .g(inst[15]));
NEMR4T g724(.s(int_128), .d(int_121), .b(gnd), .g(inst[15]));
NEMR4T g725(.s(int_129), .d(int_190), .b(gnd), .g(irq));
NEMR4T g726(.s(int_129), .d(int_123), .b(gnd), .g(ireset));
NEMR4T g727(.s(write_strobe1), .d(int_129), .b(vdd), .g(clk));
NEMR4T g728(.s(write_strobe), .d(write_strobe20), .b(vdd), .g(inst[16]));
NEMR4T g729(.s(write_strobe20), .d(int_221), .b(gnd), .g(clk));
NEMR4T g730(.s(next_interrupt_enabled), .d(next_interrupt_enabled0), .b(vdd), .g(interrupt_enabled));
NEMR4T g731(.s(next_interrupt_enabled0), .d(next_interrupt_enabled00), .b(vdd), .g(inst[13]));
NEMR4T g732(.s(next_interrupt_enabled00), .d(int_223), .b(vdd), .g(inst[16]));
NEMR4T g733(.s(int_223), .d(int_193), .b(vdd), .g(irq));
NEMR4T g734(.s(int_193), .d(int_130), .b(vdd), .g(ireset));
NEMR4T g735(.s(int_130), .d(int_13), .b(gnd), .g(inst[15]));
NEMR4T g736(.s(next_interrupt_enabled00), .d(next_interrupt_enabled001), .b(gnd), .g(inst[16]));
NEMR4T g737(.s(next_interrupt_enabled001), .d(int_39), .b(vdd), .g(irq));
NEMR4T g738(.s(next_interrupt_enabled001), .d(int_92), .b(gnd), .g(irq));
NEMR4T g739(.s(next_interrupt_enabled0), .d(int_223), .b(gnd), .g(inst[13]));
NEMR4T g740(.s(next_interrupt_enabled0), .d(int_154), .b(vdd), .g(irq));
NEMR4T g741(.s(next_interrupt_enabled), .d(next_interrupt_enabled1), .b(gnd), .g(interrupt_enabled));
NEMR4T g742(.s(next_interrupt_enabled1), .d(next_interrupt_enabled10), .b(vdd), .g(inst[13]));
NEMR4T g743(.s(next_interrupt_enabled10), .d(int_180), .b(vdd), .g(inst[16]));
NEMR4T g744(.s(next_interrupt_enabled10), .d(int_92), .b(gnd), .g(inst[16]));
NEMR4T g745(.s(next_interrupt_enabled1), .d(int_180), .b(gnd), .g(inst[13]));
NEMR4T g746(.s(next_interrupt_enabled1), .d(next_interrupt_enabled12220), .b(vdd), .g(irq));
NEMR4T g747(.s(next_interrupt_enabled12220), .d(next_interrupt_enabled122200), .b(vdd), .g(ireset));
NEMR4T g748(.s(next_interrupt_enabled122200), .d(int_0), .b(vdd), .g(inst[15]));
NEMR4T g749(.s(next_interrupt_enabled122200), .d(int_15), .b(gnd), .g(inst[15]));
NEMR4T g750(.s(next_interrupt_enabled), .d(next_interrupt_enabled20), .b(vdd), .g(inst[13]));
NEMR4T g751(.s(next_interrupt_enabled20), .d(int_92), .b(vdd), .g(inst[16]));
NEMR4T g752(.s(next_interrupt_enabled20), .d(next_interrupt_enabled201), .b(gnd), .g(inst[16]));
NEMR4T g753(.s(next_interrupt_enabled201), .d(int_93), .b(vdd), .g(inst[0]));
NEMR4T g754(.s(next_interrupt_enabled201), .d(int_180), .b(gnd), .g(inst[0]));
NEMR4T g755(.s(next_interrupt_enabled), .d(int_92), .b(gnd), .g(inst[13]));
NEMR4T g756(.s(next_interrupt_enabled), .d(int_145), .b(gnd), .g(irq));
NEMR4T g757(.s(next_interrupt_enabled), .d(int_99), .b(gnd), .g(ireset));
NEMR4T g758(.s(werf), .d(werf0), .b(vdd), .g(inst[17]));
NEMR4T g759(.s(werf0), .d(werf00), .b(vdd), .g(irq));
NEMR4T g760(.s(werf00), .d(werf000), .b(vdd), .g(ireset));
NEMR4T g761(.s(werf000), .d(werf0001), .b(gnd), .g(inst[15]));
NEMR4T g762(.s(werf0001), .d(werf00010), .b(vdd), .g(inst[14]));
NEMR4T g763(.s(werf00010), .d(int_131), .b(gnd), .g(inst[13]));
NEMR4T g764(.s(int_131), .d(vdd), .b(vdd), .g(inst[16]));
NEMR4T g765(.s(werf0001), .d(vdd), .b(gnd), .g(inst[16]));
NEMR4T g766(.s(werf000), .d(int_131), .b(gnd), .g(inst[14]));
NEMR4T g767(.s(werf0), .d(werf01), .b(gnd), .g(irq));
NEMR4T g768(.s(werf01), .d(werf011), .b(gnd), .g(ireset));
NEMR4T g769(.s(werf011), .d(int_224), .b(gnd), .g(inst[15]));
NEMR4T g770(.s(int_224), .d(int_194), .b(vdd), .g(inst[14]));
NEMR4T g771(.s(int_194), .d(int_132), .b(vdd), .g(inst[13]));
NEMR4T g772(.s(int_132), .d(gnd), .b(vdd), .g(inst[16]));
NEMR4T g773(.s(werf0), .d(werf021), .b(gnd), .g(ireset));
NEMR4T g774(.s(werf021), .d(int_134), .b(gnd), .g(inst[15]));
NEMR4T g775(.s(int_134), .d(int_133), .b(vdd), .g(inst[14]));
NEMR4T g776(.s(int_133), .d(int_132), .b(gnd), .g(inst[13]));
NEMR4T g777(.s(int_134), .d(int_132), .b(gnd), .g(inst[14]));
NEMR4T g778(.s(int_134), .d(gnd), .b(gnd), .g(inst[16]));
NEMR4T g779(.s(werf), .d(werf1), .b(gnd), .g(inst[17]));
NEMR4T g780(.s(werf1), .d(werf10), .b(vdd), .g(irq));
NEMR4T g781(.s(werf10), .d(werf100), .b(vdd), .g(ireset));
NEMR4T g782(.s(werf100), .d(werf1000), .b(vdd), .g(inst[15]));
NEMR4T g783(.s(werf1000), .d(int_132), .b(gnd), .g(inst[14]));
NEMR4T g784(.s(werf10), .d(int_134), .b(gnd), .g(inst[15]));
NEMR4T g785(.s(werf1), .d(werf11), .b(gnd), .g(irq));
NEMR4T g786(.s(werf11), .d(int_130), .b(gnd), .g(ireset));
NEMR4T g787(.s(werf), .d(werf20), .b(vdd), .g(irq));
NEMR4T g788(.s(werf20), .d(werf200), .b(vdd), .g(ireset));
NEMR4T g789(.s(werf200), .d(werf2000), .b(vdd), .g(inst[15]));
NEMR4T g790(.s(werf2000), .d(werf20000), .b(vdd), .g(inst[14]));
NEMR4T g791(.s(werf20000), .d(werf200000), .b(vdd), .g(inst[13]));
NEMR4T g792(.s(werf200000), .d(vdd), .b(vdd), .g(inst[16]));
NEMR4T g793(.s(werf200000), .d(gnd), .b(gnd), .g(inst[16]));
NEMR4T g794(.s(werf20000), .d(int_13), .b(gnd), .g(inst[13]));
NEMR4T g795(.s(werf2000), .d(werf20001), .b(gnd), .g(inst[14]));
NEMR4T g796(.s(werf20001), .d(gnd), .b(gnd), .g(inst[16]));
NEMR4T g797(.s(werf20), .d(int_224), .b(gnd), .g(inst[15]));
NEMR4T g798(.s(werf), .d(int_145), .b(gnd), .g(irq));
NEMR4T g799(.s(werf), .d(int_36), .b(gnd), .g(ireset));
NEMR4T g800(.s(wesp), .d(wesp0), .b(vdd), .g(irq));
NEMR4T g801(.s(wesp0), .d(wesp00), .b(vdd), .g(ireset));
NEMR4T g802(.s(wesp00), .d(int_196), .b(vdd), .g(inst[15]));
NEMR4T g803(.s(int_196), .d(int_195), .b(vdd), .g(inst[16]));
NEMR4T g804(.s(int_195), .d(int_135), .b(vdd), .g(inst[14]));
NEMR4T g805(.s(int_135), .d(gnd), .b(vdd), .g(inst[13]));
NEMR4T g806(.s(int_196), .d(int_135), .b(gnd), .g(inst[16]));
NEMR4T g807(.s(int_196), .d(gnd), .b(gnd), .g(inst[13]));
NEMR4T g808(.s(wesp00), .d(wesp001), .b(gnd), .g(inst[15]));
NEMR4T g809(.s(wesp001), .d(wesp0011), .b(gnd), .g(inst[17]));
NEMR4T g810(.s(wesp0011), .d(wesp00110), .b(vdd), .g(inst[16]));
NEMR4T g811(.s(wesp00110), .d(int_13), .b(vdd), .g(inst[14]));
NEMR4T g812(.s(wesp00110), .d(wesp001101), .b(gnd), .g(inst[14]));
NEMR4T g813(.s(wesp001101), .d(vdd), .b(gnd), .g(inst[13]));
NEMR4T g814(.s(wesp0011), .d(int_13), .b(gnd), .g(inst[16]));
NEMR4T g815(.s(wesp0), .d(wesp01), .b(gnd), .g(ireset));
NEMR4T g816(.s(wesp01), .d(wesp011), .b(gnd), .g(inst[15]));
NEMR4T g817(.s(wesp011), .d(int_197), .b(vdd), .g(inst[17]));
NEMR4T g818(.s(int_197), .d(int_136), .b(vdd), .g(inst[16]));
NEMR4T g819(.s(int_136), .d(int_135), .b(gnd), .g(inst[14]));
NEMR4T g820(.s(wesp0), .d(wesp021), .b(gnd), .g(inst[15]));
NEMR4T g821(.s(wesp021), .d(int_196), .b(vdd), .g(inst[17]));
NEMR4T g822(.s(wesp), .d(wesp1), .b(gnd), .g(irq));
NEMR4T g823(.s(wesp1), .d(int_196), .b(vdd), .g(ireset));
NEMR4T g824(.s(wesp1), .d(int_122), .b(gnd), .g(ireset));
NEMR4T g825(.s(wesp), .d(int_197), .b(vdd), .g(ireset));
NEMR4T g826(.s(wesp), .d(int_123), .b(gnd), .g(ireset));

endmodule
