module Instruction_decode(clk, ireset, irq, inst, c, z, read_strobe,
     write_strobe, interrupt_ack, next_interrupt_enabled,
     interrupt_enabled, zsel, csel, wsel, pcsel, stsel, werf, wesp);
  input clk, ireset, irq, c, z, interrupt_enabled;
  input [17:0] inst;
  output read_strobe, write_strobe, interrupt_ack,
       next_interrupt_enabled, werf, wesp;
  output [2:0] zsel, csel, wsel;
  output [1:0] pcsel, stsel;

  wire AA_100, AA_101, AA_102, AA_104, AA_105, AA_106, AA_107, AA_108, AA_128, AA_132, 
       AA_157, AA_158, AA_159, AA_160, AA_165, AA_166, AA_169, AA_170, AA_171, AA_172, 
       AA_173, AA_174, AA_178, AA_182, AA_200, AA_201, AA_207, AA_208, AA_210, AA_211, 
       AA_212, AA_213, AA_217, AA_218, AA_219, AA_220, AA_221, AA_222, AA_223, AA_224, 
       AA_225, AA_236, AA_244, AA_245, AA_246, AA_247, AA_248, AA_250, AA_251, AA_254, 
       AA_255, AA_256, AA_257, AA_258, AA_265, AA_283, AA_284, AA_285, AA_289, AA_290, 
       AA_291, AA_292, AA_293, AA_315, AA_316, AA_344, AA_345, AA_360, AA_361, AA_362, 
       AA_374, AA_375, AA_378, AA_379, AA_382, AA_385, AA_386, AA_387, AA_388, AA_394, 
       AA_395, AA_396, AA_397, AA_398, AA_399, AA_40, AA_400, AA_401, AA_402, AA_403, 
       AA_404, AA_49, AA_50, AA_51, AA_53, AA_84, AA_85, AA_86, AA_89, AA_99, 
       csel[0], csel[0]0, csel[0]00, csel[0]1, csel[0]10, csel[1], csel[1]0, csel[1]00, csel[1]1, csel[1]10, 
       csel[2], csel[2]0, csel[2]00, csel[2]01, interrupt_ack, interrupt_ack0, interrupt_ack1, next_interrupt_enabled, next_interrupt_enabled0, next_interrupt_enabled1, 
       next_interrupt_enabled10, next_interrupt_enabled101, next_interrupt_enabled1010, next_interrupt_enabled10100, next_interrupt_enabled11, pcsel[0], pcsel[0]0, pcsel[0]1, pcsel[0]10, pcsel[0]100, 
       pcsel[0]101, pcsel[0]11, pcsel[0]110, pcsel[0]111, pcsel[1], pcsel[1]0, pcsel[1]1, pcsel[1]10, pcsel[1]100, pcsel[1]101, 
       pcsel[1]11, pcsel[1]110, pcsel[1]111, read_strobe, read_strobe1, read_strobe10, stsel[0], stsel[0]0, stsel[0]1, stsel[0]10, 
       stsel[0]100, stsel[0]101, stsel[0]11, stsel[0]110, stsel[0]111, stsel[1], stsel[1]0, stsel[1]1, stsel[1]10, stsel[1]100, 
       stsel[1]101, stsel[1]11, stsel[1]110, stsel[1]111, werf, werf0, werf00, werf000, werf0000, werf1, 
       werf10, wesp, wesp1, write_strobe, write_strobe0, write_strobe01, write_strobe1, wsel[0], wsel[0]0, wsel[0]1, 
       wsel[0]10, wsel[1], zsel[0], zsel[0]0, zsel[0]00, zsel[0]1, zsel[0]11, zsel[0]110, zsel[0]1100, zsel[1], 
       zsel[1]0, zsel[1]00, zsel[1]01, zsel[1]1, zsel[2], zsel[2]0, zsel[2]1;

assign wsel[2] = inst[16];

NEMR4T g1(.s(zsel[0]), .d(zsel[0]0), .b(vdd), .g(inst[14]));
NEMR4T g2(.s(zsel[0]0), .d(zsel[0]00), .b(vdd), .g(inst[16]));
NEMR4T g3(.s(zsel[0]00), .d(AA_107), .b(vdd), .g(inst[13]));
NEMR4T g4(.s(AA_107), .d(AA_221), .b(vdd), .g(irq));
NEMR4T g5(.s(AA_221), .d(AA_220), .b(vdd), .g(inst[17]));
NEMR4T g6(.s(AA_220), .d(AA_394), .b(vdd), .g(ireset));
NEMR4T g7(.s(AA_394), .d(gnd), .b(vdd), .g(inst[15]));
NEMR4T g8(.s(AA_394), .d(gnd), .b(gnd), .g(inst[15]));
NEMR4T g9(.s(AA_220), .d(AA_378), .b(gnd), .g(ireset));
NEMR4T g10(.s(AA_378), .d(vdd), .b(vdd), .g(inst[15]));
NEMR4T g11(.s(AA_378), .d(vdd), .b(gnd), .g(inst[15]));
NEMR4T g12(.s(AA_221), .d(AA_217), .b(gnd), .g(inst[17]));
NEMR4T g13(.s(AA_217), .d(AA_379), .b(vdd), .g(ireset));
NEMR4T g14(.s(AA_379), .d(vdd), .b(vdd), .g(inst[15]));
NEMR4T g15(.s(AA_379), .d(gnd), .b(gnd), .g(inst[15]));
NEMR4T g16(.s(AA_217), .d(AA_378), .b(gnd), .g(ireset));
NEMR4T g17(.s(AA_107), .d(AA_222), .b(gnd), .g(irq));
NEMR4T g18(.s(AA_222), .d(AA_220), .b(vdd), .g(inst[17]));
NEMR4T g19(.s(AA_222), .d(AA_220), .b(gnd), .g(inst[17]));
NEMR4T g20(.s(zsel[0]00), .d(AA_99), .b(gnd), .g(inst[13]));
NEMR4T g21(.s(AA_99), .d(AA_222), .b(vdd), .g(irq));
NEMR4T g22(.s(AA_99), .d(AA_222), .b(gnd), .g(irq));
NEMR4T g23(.s(zsel[0]0), .d(AA_102), .b(gnd), .g(inst[16]));
NEMR4T g24(.s(AA_102), .d(AA_101), .b(vdd), .g(inst[13]));
NEMR4T g25(.s(AA_101), .d(AA_100), .b(vdd), .g(irq));
NEMR4T g26(.s(AA_100), .d(AA_178), .b(vdd), .g(inst[17]));
NEMR4T g27(.s(AA_178), .d(AA_395), .b(vdd), .g(ireset));
NEMR4T g28(.s(AA_395), .d(gnd), .b(vdd), .g(inst[15]));
NEMR4T g29(.s(AA_395), .d(vdd), .b(gnd), .g(inst[15]));
NEMR4T g30(.s(AA_178), .d(AA_378), .b(gnd), .g(ireset));
NEMR4T g31(.s(AA_100), .d(AA_220), .b(gnd), .g(inst[17]));
NEMR4T g32(.s(AA_101), .d(AA_222), .b(gnd), .g(irq));
NEMR4T g33(.s(AA_102), .d(AA_101), .b(gnd), .g(inst[13]));
NEMR4T g34(.s(zsel[0]), .d(zsel[0]1), .b(gnd), .g(inst[14]));
NEMR4T g35(.s(zsel[0]1), .d(AA_40), .b(vdd), .g(inst[16]));
NEMR4T g36(.s(AA_40), .d(AA_99), .b(vdd), .g(inst[13]));
NEMR4T g37(.s(AA_40), .d(AA_99), .b(gnd), .g(inst[13]));
NEMR4T g38(.s(zsel[0]1), .d(zsel[0]11), .b(gnd), .g(inst[16]));
NEMR4T g39(.s(zsel[0]11), .d(zsel[0]110), .b(vdd), .g(inst[13]));
NEMR4T g40(.s(zsel[0]110), .d(zsel[0]1100), .b(vdd), .g(irq));
NEMR4T g41(.s(zsel[0]1100), .d(AA_218), .b(vdd), .g(inst[17]));
NEMR4T g42(.s(AA_218), .d(AA_378), .b(vdd), .g(ireset));
NEMR4T g43(.s(AA_218), .d(AA_378), .b(gnd), .g(ireset));
NEMR4T g44(.s(zsel[0]1100), .d(AA_220), .b(gnd), .g(inst[17]));
NEMR4T g45(.s(zsel[0]110), .d(AA_222), .b(gnd), .g(irq));
NEMR4T g46(.s(zsel[0]11), .d(AA_101), .b(gnd), .g(inst[13]));
NEMR4T g47(.s(zsel[1]), .d(zsel[1]0), .b(vdd), .g(inst[14]));
NEMR4T g48(.s(zsel[1]0), .d(zsel[1]00), .b(vdd), .g(inst[16]));
NEMR4T g49(.s(zsel[1]00), .d(AA_128), .b(vdd), .g(inst[13]));
NEMR4T g50(.s(AA_128), .d(AA_265), .b(vdd), .g(irq));
NEMR4T g51(.s(AA_265), .d(AA_396), .b(vdd), .g(inst[17]));
NEMR4T g52(.s(AA_396), .d(AA_394), .b(vdd), .g(ireset));
NEMR4T g53(.s(AA_396), .d(AA_394), .b(gnd), .g(ireset));
NEMR4T g54(.s(AA_265), .d(AA_382), .b(gnd), .g(inst[17]));
NEMR4T g55(.s(AA_382), .d(AA_379), .b(vdd), .g(ireset));
NEMR4T g56(.s(AA_382), .d(AA_394), .b(gnd), .g(ireset));
NEMR4T g57(.s(AA_128), .d(AA_397), .b(gnd), .g(irq));
NEMR4T g58(.s(AA_397), .d(AA_396), .b(vdd), .g(inst[17]));
NEMR4T g59(.s(AA_397), .d(AA_396), .b(gnd), .g(inst[17]));
NEMR4T g60(.s(zsel[1]00), .d(AA_386), .b(gnd), .g(inst[13]));
NEMR4T g61(.s(AA_386), .d(AA_385), .b(vdd), .g(irq));
NEMR4T g62(.s(AA_385), .d(AA_398), .b(vdd), .g(inst[17]));
NEMR4T g63(.s(AA_398), .d(AA_395), .b(vdd), .g(ireset));
NEMR4T g64(.s(AA_398), .d(AA_394), .b(gnd), .g(ireset));
NEMR4T g65(.s(AA_385), .d(AA_396), .b(gnd), .g(inst[17]));
NEMR4T g66(.s(AA_386), .d(AA_397), .b(gnd), .g(irq));
NEMR4T g67(.s(zsel[1]0), .d(zsel[1]01), .b(gnd), .g(inst[16]));
NEMR4T g68(.s(zsel[1]01), .d(AA_399), .b(vdd), .g(inst[13]));
NEMR4T g69(.s(AA_399), .d(AA_397), .b(vdd), .g(irq));
NEMR4T g70(.s(AA_399), .d(AA_397), .b(gnd), .g(irq));
NEMR4T g71(.s(zsel[1]01), .d(AA_316), .b(gnd), .g(inst[13]));
NEMR4T g72(.s(AA_316), .d(AA_315), .b(vdd), .g(irq));
NEMR4T g73(.s(AA_315), .d(AA_382), .b(vdd), .g(inst[17]));
NEMR4T g74(.s(AA_315), .d(AA_396), .b(gnd), .g(inst[17]));
NEMR4T g75(.s(AA_316), .d(AA_397), .b(gnd), .g(irq));
NEMR4T g76(.s(zsel[1]), .d(zsel[1]1), .b(gnd), .g(inst[14]));
NEMR4T g77(.s(zsel[1]1), .d(AA_387), .b(vdd), .g(inst[16]));
NEMR4T g78(.s(AA_387), .d(AA_386), .b(vdd), .g(inst[13]));
NEMR4T g79(.s(AA_387), .d(AA_386), .b(gnd), .g(inst[13]));
NEMR4T g80(.s(zsel[1]1), .d(AA_400), .b(gnd), .g(inst[16]));
NEMR4T g81(.s(AA_400), .d(AA_399), .b(vdd), .g(inst[13]));
NEMR4T g82(.s(AA_400), .d(AA_399), .b(gnd), .g(inst[13]));
NEMR4T g83(.s(zsel[2]), .d(zsel[2]0), .b(vdd), .g(inst[14]));
NEMR4T g84(.s(zsel[2]0), .d(AA_40), .b(vdd), .g(inst[16]));
NEMR4T g85(.s(zsel[2]0), .d(AA_105), .b(gnd), .g(inst[16]));
NEMR4T g86(.s(AA_105), .d(AA_104), .b(vdd), .g(inst[13]));
NEMR4T g87(.s(AA_104), .d(AA_182), .b(vdd), .g(irq));
NEMR4T g88(.s(AA_182), .d(AA_220), .b(vdd), .g(inst[17]));
NEMR4T g89(.s(AA_182), .d(AA_178), .b(gnd), .g(inst[17]));
NEMR4T g90(.s(AA_104), .d(AA_222), .b(gnd), .g(irq));
NEMR4T g91(.s(AA_105), .d(AA_99), .b(gnd), .g(inst[13]));
NEMR4T g92(.s(zsel[2]), .d(zsel[2]1), .b(gnd), .g(inst[14]));
NEMR4T g93(.s(zsel[2]1), .d(AA_40), .b(vdd), .g(inst[16]));
NEMR4T g94(.s(zsel[2]1), .d(AA_40), .b(gnd), .g(inst[16]));
NEMR4T g95(.s(csel[0]), .d(csel[0]0), .b(vdd), .g(inst[3]));
NEMR4T g96(.s(csel[0]0), .d(csel[0]00), .b(vdd), .g(inst[14]));
NEMR4T g97(.s(csel[0]00), .d(AA_106), .b(vdd), .g(inst[16]));
NEMR4T g98(.s(AA_106), .d(AA_99), .b(vdd), .g(inst[13]));
NEMR4T g99(.s(AA_106), .d(AA_101), .b(gnd), .g(inst[13]));
NEMR4T g100(.s(csel[0]00), .d(AA_51), .b(gnd), .g(inst[16]));
NEMR4T g101(.s(AA_51), .d(AA_50), .b(vdd), .g(inst[13]));
NEMR4T g102(.s(AA_50), .d(AA_49), .b(vdd), .g(irq));
NEMR4T g103(.s(AA_49), .d(AA_178), .b(vdd), .g(inst[17]));
NEMR4T g104(.s(AA_49), .d(AA_178), .b(gnd), .g(inst[17]));
NEMR4T g105(.s(AA_50), .d(AA_222), .b(gnd), .g(irq));
NEMR4T g106(.s(AA_51), .d(AA_101), .b(gnd), .g(inst[13]));
NEMR4T g107(.s(csel[0]0), .d(AA_53), .b(gnd), .g(inst[14]));
NEMR4T g108(.s(AA_53), .d(AA_102), .b(vdd), .g(inst[16]));
NEMR4T g109(.s(AA_53), .d(AA_102), .b(gnd), .g(inst[16]));
NEMR4T g110(.s(csel[0]), .d(csel[0]1), .b(gnd), .g(inst[3]));
NEMR4T g111(.s(csel[0]1), .d(csel[0]10), .b(vdd), .g(inst[14]));
NEMR4T g112(.s(csel[0]10), .d(AA_108), .b(vdd), .g(inst[16]));
NEMR4T g113(.s(AA_108), .d(AA_107), .b(vdd), .g(inst[13]));
NEMR4T g114(.s(AA_108), .d(AA_101), .b(gnd), .g(inst[13]));
NEMR4T g115(.s(csel[0]10), .d(AA_51), .b(gnd), .g(inst[16]));
NEMR4T g116(.s(csel[0]1), .d(AA_53), .b(gnd), .g(inst[14]));
NEMR4T g117(.s(csel[1]), .d(csel[1]0), .b(vdd), .g(inst[3]));
NEMR4T g118(.s(csel[1]0), .d(csel[1]00), .b(vdd), .g(inst[14]));
NEMR4T g119(.s(csel[1]00), .d(AA_108), .b(vdd), .g(inst[16]));
NEMR4T g120(.s(csel[1]00), .d(AA_105), .b(gnd), .g(inst[16]));
NEMR4T g121(.s(csel[1]0), .d(AA_89), .b(gnd), .g(inst[14]));
NEMR4T g122(.s(AA_89), .d(AA_102), .b(vdd), .g(inst[16]));
NEMR4T g123(.s(AA_89), .d(AA_86), .b(gnd), .g(inst[16]));
NEMR4T g124(.s(AA_86), .d(AA_85), .b(vdd), .g(inst[13]));
NEMR4T g125(.s(AA_85), .d(AA_84), .b(vdd), .g(irq));
NEMR4T g126(.s(AA_84), .d(AA_217), .b(vdd), .g(inst[17]));
NEMR4T g127(.s(AA_84), .d(AA_220), .b(gnd), .g(inst[17]));
NEMR4T g128(.s(AA_85), .d(AA_222), .b(gnd), .g(irq));
NEMR4T g129(.s(AA_86), .d(AA_99), .b(gnd), .g(inst[13]));
NEMR4T g130(.s(csel[1]), .d(csel[1]1), .b(gnd), .g(inst[3]));
NEMR4T g131(.s(csel[1]1), .d(csel[1]10), .b(vdd), .g(inst[14]));
NEMR4T g132(.s(csel[1]10), .d(AA_106), .b(vdd), .g(inst[16]));
NEMR4T g133(.s(csel[1]10), .d(AA_105), .b(gnd), .g(inst[16]));
NEMR4T g134(.s(csel[1]1), .d(AA_89), .b(gnd), .g(inst[14]));
NEMR4T g135(.s(csel[2]), .d(csel[2]0), .b(vdd), .g(inst[14]));
NEMR4T g136(.s(csel[2]0), .d(csel[2]00), .b(vdd), .g(inst[16]));
NEMR4T g137(.s(csel[2]00), .d(AA_128), .b(vdd), .g(inst[13]));
NEMR4T g138(.s(csel[2]00), .d(AA_399), .b(gnd), .g(inst[13]));
NEMR4T g139(.s(csel[2]0), .d(csel[2]01), .b(gnd), .g(inst[16]));
NEMR4T g140(.s(csel[2]01), .d(AA_402), .b(vdd), .g(inst[13]));
NEMR4T g141(.s(AA_402), .d(AA_401), .b(vdd), .g(irq));
NEMR4T g142(.s(AA_401), .d(AA_396), .b(vdd), .g(inst[17]));
NEMR4T g143(.s(AA_401), .d(AA_398), .b(gnd), .g(inst[17]));
NEMR4T g144(.s(AA_402), .d(AA_397), .b(gnd), .g(irq));
NEMR4T g145(.s(csel[2]01), .d(AA_316), .b(gnd), .g(inst[13]));
NEMR4T g146(.s(csel[2]), .d(AA_403), .b(gnd), .g(inst[14]));
NEMR4T g147(.s(AA_403), .d(AA_400), .b(vdd), .g(inst[16]));
NEMR4T g148(.s(AA_403), .d(AA_400), .b(gnd), .g(inst[16]));
NEMR4T g149(.s(wsel[0]), .d(wsel[0]0), .b(vdd), .g(inst[14]));
NEMR4T g150(.s(wsel[0]0), .d(AA_132), .b(vdd), .g(inst[13]));
NEMR4T g151(.s(AA_132), .d(AA_394), .b(vdd), .g(inst[17]));
NEMR4T g152(.s(AA_132), .d(AA_378), .b(gnd), .g(inst[17]));
NEMR4T g153(.s(wsel[0]0), .d(AA_132), .b(gnd), .g(inst[13]));
NEMR4T g154(.s(wsel[0]), .d(wsel[0]1), .b(gnd), .g(inst[14]));
NEMR4T g155(.s(wsel[0]1), .d(wsel[0]10), .b(vdd), .g(inst[13]));
NEMR4T g156(.s(wsel[0]10), .d(AA_379), .b(vdd), .g(inst[17]));
NEMR4T g157(.s(wsel[0]10), .d(AA_378), .b(gnd), .g(inst[17]));
NEMR4T g158(.s(wsel[0]1), .d(AA_132), .b(gnd), .g(inst[13]));
NEMR4T g159(.s(wsel[1]), .d(AA_394), .b(vdd), .g(inst[14]));
NEMR4T g160(.s(wsel[1]), .d(AA_379), .b(gnd), .g(inst[14]));
NEMR4T g161(.s(pcsel[1]), .d(pcsel[1]0), .b(vdd), .g(inst[12]));
NEMR4T g162(.s(pcsel[1]0), .d(AA_174), .b(vdd), .g(z));
NEMR4T g163(.s(AA_174), .d(AA_173), .b(vdd), .g(c));
NEMR4T g164(.s(AA_173), .d(AA_172), .b(vdd), .g(inst[11]));
NEMR4T g165(.s(AA_172), .d(AA_171), .b(vdd), .g(inst[10]));
NEMR4T g166(.s(AA_171), .d(AA_170), .b(vdd), .g(inst[14]));
NEMR4T g167(.s(AA_170), .d(AA_169), .b(vdd), .g(inst[16]));
NEMR4T g168(.s(AA_169), .d(AA_223), .b(vdd), .g(inst[13]));
NEMR4T g169(.s(AA_223), .d(AA_222), .b(vdd), .g(irq));
NEMR4T g170(.s(AA_223), .d(AA_219), .b(gnd), .g(irq));
NEMR4T g171(.s(AA_219), .d(AA_218), .b(vdd), .g(inst[17]));
NEMR4T g172(.s(AA_219), .d(AA_218), .b(gnd), .g(inst[17]));
NEMR4T g173(.s(AA_169), .d(AA_165), .b(gnd), .g(inst[13]));
NEMR4T g174(.s(AA_165), .d(AA_182), .b(vdd), .g(irq));
NEMR4T g175(.s(AA_165), .d(AA_219), .b(gnd), .g(irq));
NEMR4T g176(.s(AA_170), .d(AA_166), .b(gnd), .g(inst[16]));
NEMR4T g177(.s(AA_166), .d(AA_165), .b(vdd), .g(inst[13]));
NEMR4T g178(.s(AA_166), .d(AA_223), .b(gnd), .g(inst[13]));
NEMR4T g179(.s(AA_171), .d(AA_225), .b(gnd), .g(inst[14]));
NEMR4T g180(.s(AA_225), .d(AA_224), .b(vdd), .g(inst[16]));
NEMR4T g181(.s(AA_224), .d(AA_223), .b(vdd), .g(inst[13]));
NEMR4T g182(.s(AA_224), .d(AA_223), .b(gnd), .g(inst[13]));
NEMR4T g183(.s(AA_225), .d(AA_224), .b(gnd), .g(inst[16]));
NEMR4T g184(.s(AA_172), .d(AA_171), .b(gnd), .g(inst[10]));
NEMR4T g185(.s(AA_173), .d(AA_172), .b(gnd), .g(inst[11]));
NEMR4T g186(.s(AA_174), .d(AA_173), .b(gnd), .g(c));
NEMR4T g187(.s(pcsel[1]0), .d(AA_174), .b(gnd), .g(z));
NEMR4T g188(.s(pcsel[1]), .d(pcsel[1]1), .b(gnd), .g(inst[12]));
NEMR4T g189(.s(pcsel[1]1), .d(pcsel[1]10), .b(vdd), .g(z));
NEMR4T g190(.s(pcsel[1]10), .d(pcsel[1]100), .b(vdd), .g(c));
NEMR4T g191(.s(pcsel[1]100), .d(AA_159), .b(vdd), .g(inst[11]));
NEMR4T g192(.s(AA_159), .d(AA_158), .b(vdd), .g(inst[10]));
NEMR4T g193(.s(AA_158), .d(AA_157), .b(vdd), .g(inst[14]));
NEMR4T g194(.s(AA_157), .d(AA_224), .b(vdd), .g(inst[16]));
NEMR4T g195(.s(AA_157), .d(AA_166), .b(gnd), .g(inst[16]));
NEMR4T g196(.s(AA_158), .d(AA_225), .b(gnd), .g(inst[14]));
NEMR4T g197(.s(AA_159), .d(AA_171), .b(gnd), .g(inst[10]));
NEMR4T g198(.s(pcsel[1]100), .d(AA_159), .b(gnd), .g(inst[11]));
NEMR4T g199(.s(pcsel[1]10), .d(pcsel[1]101), .b(gnd), .g(c));
NEMR4T g200(.s(pcsel[1]101), .d(AA_159), .b(vdd), .g(inst[11]));
NEMR4T g201(.s(pcsel[1]101), .d(AA_160), .b(gnd), .g(inst[11]));
NEMR4T g202(.s(AA_160), .d(AA_171), .b(vdd), .g(inst[10]));
NEMR4T g203(.s(AA_160), .d(AA_158), .b(gnd), .g(inst[10]));
NEMR4T g204(.s(pcsel[1]1), .d(pcsel[1]11), .b(gnd), .g(z));
NEMR4T g205(.s(pcsel[1]11), .d(pcsel[1]110), .b(vdd), .g(c));
NEMR4T g206(.s(pcsel[1]110), .d(AA_160), .b(vdd), .g(inst[11]));
NEMR4T g207(.s(pcsel[1]110), .d(AA_159), .b(gnd), .g(inst[11]));
NEMR4T g208(.s(pcsel[1]11), .d(pcsel[1]111), .b(gnd), .g(c));
NEMR4T g209(.s(pcsel[1]111), .d(AA_160), .b(vdd), .g(inst[11]));
NEMR4T g210(.s(pcsel[1]111), .d(AA_160), .b(gnd), .g(inst[11]));
NEMR4T g211(.s(pcsel[0]), .d(pcsel[0]0), .b(vdd), .g(inst[12]));
NEMR4T g212(.s(pcsel[0]0), .d(AA_213), .b(vdd), .g(z));
NEMR4T g213(.s(AA_213), .d(AA_212), .b(vdd), .g(c));
NEMR4T g214(.s(AA_212), .d(AA_211), .b(vdd), .g(inst[11]));
NEMR4T g215(.s(AA_211), .d(AA_210), .b(vdd), .g(inst[10]));
NEMR4T g216(.s(AA_210), .d(AA_224), .b(vdd), .g(inst[16]));
NEMR4T g217(.s(AA_210), .d(AA_208), .b(gnd), .g(inst[16]));
NEMR4T g218(.s(AA_208), .d(AA_207), .b(vdd), .g(inst[13]));
NEMR4T g219(.s(AA_207), .d(AA_221), .b(vdd), .g(irq));
NEMR4T g220(.s(AA_207), .d(AA_219), .b(gnd), .g(irq));
NEMR4T g221(.s(AA_208), .d(AA_223), .b(gnd), .g(inst[13]));
NEMR4T g222(.s(AA_211), .d(AA_210), .b(gnd), .g(inst[10]));
NEMR4T g223(.s(AA_212), .d(AA_211), .b(gnd), .g(inst[11]));
NEMR4T g224(.s(AA_213), .d(AA_212), .b(gnd), .g(c));
NEMR4T g225(.s(pcsel[0]0), .d(AA_213), .b(gnd), .g(z));
NEMR4T g226(.s(pcsel[0]), .d(pcsel[0]1), .b(gnd), .g(inst[12]));
NEMR4T g227(.s(pcsel[0]1), .d(pcsel[0]10), .b(vdd), .g(z));
NEMR4T g228(.s(pcsel[0]10), .d(pcsel[0]100), .b(vdd), .g(c));
NEMR4T g229(.s(pcsel[0]100), .d(AA_200), .b(vdd), .g(inst[11]));
NEMR4T g230(.s(AA_200), .d(AA_225), .b(vdd), .g(inst[10]));
NEMR4T g231(.s(AA_200), .d(AA_210), .b(gnd), .g(inst[10]));
NEMR4T g232(.s(pcsel[0]100), .d(AA_200), .b(gnd), .g(inst[11]));
NEMR4T g233(.s(pcsel[0]10), .d(pcsel[0]101), .b(gnd), .g(c));
NEMR4T g234(.s(pcsel[0]101), .d(AA_200), .b(vdd), .g(inst[11]));
NEMR4T g235(.s(pcsel[0]101), .d(AA_201), .b(gnd), .g(inst[11]));
NEMR4T g236(.s(AA_201), .d(AA_210), .b(vdd), .g(inst[10]));
NEMR4T g237(.s(AA_201), .d(AA_225), .b(gnd), .g(inst[10]));
NEMR4T g238(.s(pcsel[0]1), .d(pcsel[0]11), .b(gnd), .g(z));
NEMR4T g239(.s(pcsel[0]11), .d(pcsel[0]110), .b(vdd), .g(c));
NEMR4T g240(.s(pcsel[0]110), .d(AA_201), .b(vdd), .g(inst[11]));
NEMR4T g241(.s(pcsel[0]110), .d(AA_200), .b(gnd), .g(inst[11]));
NEMR4T g242(.s(pcsel[0]11), .d(pcsel[0]111), .b(gnd), .g(c));
NEMR4T g243(.s(pcsel[0]111), .d(AA_201), .b(vdd), .g(inst[11]));
NEMR4T g244(.s(pcsel[0]111), .d(AA_201), .b(gnd), .g(inst[11]));
NEMR4T g245(.s(stsel[0]), .d(stsel[0]0), .b(vdd), .g(inst[12]));
NEMR4T g246(.s(stsel[0]0), .d(AA_258), .b(vdd), .g(z));
NEMR4T g247(.s(AA_258), .d(AA_257), .b(vdd), .g(c));
NEMR4T g248(.s(AA_257), .d(AA_256), .b(vdd), .g(inst[11]));
NEMR4T g249(.s(AA_256), .d(AA_255), .b(vdd), .g(inst[10]));
NEMR4T g250(.s(AA_255), .d(AA_254), .b(vdd), .g(inst[14]));
NEMR4T g251(.s(AA_254), .d(AA_248), .b(vdd), .g(inst[16]));
NEMR4T g252(.s(AA_248), .d(AA_247), .b(vdd), .g(inst[13]));
NEMR4T g253(.s(AA_247), .d(AA_397), .b(vdd), .g(irq));
NEMR4T g254(.s(AA_247), .d(AA_360), .b(gnd), .g(irq));
NEMR4T g255(.s(AA_360), .d(AA_388), .b(vdd), .g(inst[17]));
NEMR4T g256(.s(AA_388), .d(AA_378), .b(vdd), .g(ireset));
NEMR4T g257(.s(AA_388), .d(AA_394), .b(gnd), .g(ireset));
NEMR4T g258(.s(AA_360), .d(AA_388), .b(gnd), .g(inst[17]));
NEMR4T g259(.s(AA_248), .d(AA_247), .b(gnd), .g(inst[13]));
NEMR4T g260(.s(AA_254), .d(AA_251), .b(gnd), .g(inst[16]));
NEMR4T g261(.s(AA_251), .d(AA_250), .b(vdd), .g(inst[13]));
NEMR4T g262(.s(AA_250), .d(AA_265), .b(vdd), .g(irq));
NEMR4T g263(.s(AA_250), .d(AA_360), .b(gnd), .g(irq));
NEMR4T g264(.s(AA_251), .d(AA_247), .b(gnd), .g(inst[13]));
NEMR4T g265(.s(AA_255), .d(AA_236), .b(gnd), .g(inst[14]));
NEMR4T g266(.s(AA_236), .d(AA_248), .b(vdd), .g(inst[16]));
NEMR4T g267(.s(AA_236), .d(AA_248), .b(gnd), .g(inst[16]));
NEMR4T g268(.s(AA_256), .d(AA_255), .b(gnd), .g(inst[10]));
NEMR4T g269(.s(AA_257), .d(AA_256), .b(gnd), .g(inst[11]));
NEMR4T g270(.s(AA_258), .d(AA_257), .b(gnd), .g(c));
NEMR4T g271(.s(stsel[0]0), .d(AA_258), .b(gnd), .g(z));
NEMR4T g272(.s(stsel[0]), .d(stsel[0]1), .b(gnd), .g(inst[12]));
NEMR4T g273(.s(stsel[0]1), .d(stsel[0]10), .b(vdd), .g(z));
NEMR4T g274(.s(stsel[0]10), .d(stsel[0]100), .b(vdd), .g(c));
NEMR4T g275(.s(stsel[0]100), .d(AA_245), .b(vdd), .g(inst[11]));
NEMR4T g276(.s(AA_245), .d(AA_244), .b(vdd), .g(inst[10]));
NEMR4T g277(.s(AA_244), .d(AA_236), .b(vdd), .g(inst[14]));
NEMR4T g278(.s(AA_244), .d(AA_236), .b(gnd), .g(inst[14]));
NEMR4T g279(.s(AA_245), .d(AA_255), .b(gnd), .g(inst[10]));
NEMR4T g280(.s(stsel[0]100), .d(AA_245), .b(gnd), .g(inst[11]));
NEMR4T g281(.s(stsel[0]10), .d(stsel[0]101), .b(gnd), .g(c));
NEMR4T g282(.s(stsel[0]101), .d(AA_245), .b(vdd), .g(inst[11]));
NEMR4T g283(.s(stsel[0]101), .d(AA_246), .b(gnd), .g(inst[11]));
NEMR4T g284(.s(AA_246), .d(AA_255), .b(vdd), .g(inst[10]));
NEMR4T g285(.s(AA_246), .d(AA_244), .b(gnd), .g(inst[10]));
NEMR4T g286(.s(stsel[0]1), .d(stsel[0]11), .b(gnd), .g(z));
NEMR4T g287(.s(stsel[0]11), .d(stsel[0]110), .b(vdd), .g(c));
NEMR4T g288(.s(stsel[0]110), .d(AA_246), .b(vdd), .g(inst[11]));
NEMR4T g289(.s(stsel[0]110), .d(AA_245), .b(gnd), .g(inst[11]));
NEMR4T g290(.s(stsel[0]11), .d(stsel[0]111), .b(gnd), .g(c));
NEMR4T g291(.s(stsel[0]111), .d(AA_246), .b(vdd), .g(inst[11]));
NEMR4T g292(.s(stsel[0]111), .d(AA_246), .b(gnd), .g(inst[11]));
NEMR4T g293(.s(stsel[1]), .d(stsel[1]0), .b(vdd), .g(inst[12]));
NEMR4T g294(.s(stsel[1]0), .d(AA_293), .b(vdd), .g(z));
NEMR4T g295(.s(AA_293), .d(AA_292), .b(vdd), .g(c));
NEMR4T g296(.s(AA_292), .d(AA_291), .b(vdd), .g(inst[11]));
NEMR4T g297(.s(AA_291), .d(AA_290), .b(vdd), .g(inst[10]));
NEMR4T g298(.s(AA_290), .d(AA_289), .b(vdd), .g(inst[14]));
NEMR4T g299(.s(AA_289), .d(AA_404), .b(vdd), .g(inst[16]));
NEMR4T g300(.s(AA_404), .d(AA_399), .b(vdd), .g(inst[13]));
NEMR4T g301(.s(AA_404), .d(AA_402), .b(gnd), .g(inst[13]));
NEMR4T g302(.s(AA_289), .d(AA_361), .b(gnd), .g(inst[16]));
NEMR4T g303(.s(AA_361), .d(AA_402), .b(vdd), .g(inst[13]));
NEMR4T g304(.s(AA_361), .d(AA_399), .b(gnd), .g(inst[13]));
NEMR4T g305(.s(AA_290), .d(AA_403), .b(gnd), .g(inst[14]));
NEMR4T g306(.s(AA_291), .d(AA_290), .b(gnd), .g(inst[10]));
NEMR4T g307(.s(AA_292), .d(AA_291), .b(gnd), .g(inst[11]));
NEMR4T g308(.s(AA_293), .d(AA_292), .b(gnd), .g(c));
NEMR4T g309(.s(stsel[1]0), .d(AA_293), .b(gnd), .g(z));
NEMR4T g310(.s(stsel[1]), .d(stsel[1]1), .b(gnd), .g(inst[12]));
NEMR4T g311(.s(stsel[1]1), .d(stsel[1]10), .b(vdd), .g(z));
NEMR4T g312(.s(stsel[1]10), .d(stsel[1]100), .b(vdd), .g(c));
NEMR4T g313(.s(stsel[1]100), .d(AA_284), .b(vdd), .g(inst[11]));
NEMR4T g314(.s(AA_284), .d(AA_283), .b(vdd), .g(inst[10]));
NEMR4T g315(.s(AA_283), .d(AA_362), .b(vdd), .g(inst[14]));
NEMR4T g316(.s(AA_362), .d(AA_400), .b(vdd), .g(inst[16]));
NEMR4T g317(.s(AA_362), .d(AA_361), .b(gnd), .g(inst[16]));
NEMR4T g318(.s(AA_283), .d(AA_403), .b(gnd), .g(inst[14]));
NEMR4T g319(.s(AA_284), .d(AA_290), .b(gnd), .g(inst[10]));
NEMR4T g320(.s(stsel[1]100), .d(AA_284), .b(gnd), .g(inst[11]));
NEMR4T g321(.s(stsel[1]10), .d(stsel[1]101), .b(gnd), .g(c));
NEMR4T g322(.s(stsel[1]101), .d(AA_284), .b(vdd), .g(inst[11]));
NEMR4T g323(.s(stsel[1]101), .d(AA_285), .b(gnd), .g(inst[11]));
NEMR4T g324(.s(AA_285), .d(AA_290), .b(vdd), .g(inst[10]));
NEMR4T g325(.s(AA_285), .d(AA_283), .b(gnd), .g(inst[10]));
NEMR4T g326(.s(stsel[1]1), .d(stsel[1]11), .b(gnd), .g(z));
NEMR4T g327(.s(stsel[1]11), .d(stsel[1]110), .b(vdd), .g(c));
NEMR4T g328(.s(stsel[1]110), .d(AA_285), .b(vdd), .g(inst[11]));
NEMR4T g329(.s(stsel[1]110), .d(AA_284), .b(gnd), .g(inst[11]));
NEMR4T g330(.s(stsel[1]11), .d(stsel[1]111), .b(gnd), .g(c));
NEMR4T g331(.s(stsel[1]111), .d(AA_285), .b(vdd), .g(inst[11]));
NEMR4T g332(.s(stsel[1]111), .d(AA_285), .b(gnd), .g(inst[11]));
NEMR4T g333(.s(read_strobe), .d(AA_403), .b(vdd), .g(inst[14]));
NEMR4T g334(.s(read_strobe), .d(read_strobe1), .b(gnd), .g(inst[14]));
NEMR4T g335(.s(read_strobe1), .d(read_strobe10), .b(vdd), .g(inst[16]));
NEMR4T g336(.s(read_strobe10), .d(AA_316), .b(vdd), .g(inst[13]));
NEMR4T g337(.s(read_strobe10), .d(AA_399), .b(gnd), .g(inst[13]));
NEMR4T g338(.s(read_strobe1), .d(AA_400), .b(gnd), .g(inst[16]));
NEMR4T g339(.s(write_strobe), .d(write_strobe0), .b(vdd), .g(clk));
NEMR4T g340(.s(write_strobe0), .d(AA_403), .b(vdd), .g(inst[14]));
NEMR4T g341(.s(write_strobe0), .d(write_strobe01), .b(gnd), .g(inst[14]));
NEMR4T g342(.s(write_strobe01), .d(AA_361), .b(vdd), .g(inst[16]));
NEMR4T g343(.s(write_strobe01), .d(AA_400), .b(gnd), .g(inst[16]));
NEMR4T g344(.s(write_strobe), .d(write_strobe1), .b(gnd), .g(clk));
NEMR4T g345(.s(write_strobe1), .d(AA_403), .b(vdd), .g(inst[14]));
NEMR4T g346(.s(write_strobe1), .d(AA_403), .b(gnd), .g(inst[14]));
NEMR4T g347(.s(interrupt_ack), .d(interrupt_ack0), .b(vdd), .g(irq));
NEMR4T g348(.s(interrupt_ack0), .d(gnd), .b(vdd), .g(ireset));
NEMR4T g349(.s(interrupt_ack0), .d(gnd), .b(gnd), .g(ireset));
NEMR4T g350(.s(interrupt_ack), .d(interrupt_ack1), .b(gnd), .g(irq));
NEMR4T g351(.s(interrupt_ack1), .d(vdd), .b(vdd), .g(ireset));
NEMR4T g352(.s(interrupt_ack1), .d(gnd), .b(gnd), .g(ireset));
NEMR4T g353(.s(next_interrupt_enabled), .d(next_interrupt_enabled0), .b(vdd), .g(interrupt_enabled));
NEMR4T g354(.s(next_interrupt_enabled0), .d(AA_403), .b(vdd), .g(inst[0]));
NEMR4T g355(.s(next_interrupt_enabled0), .d(AA_362), .b(gnd), .g(inst[0]));
NEMR4T g356(.s(next_interrupt_enabled), .d(next_interrupt_enabled1), .b(gnd), .g(interrupt_enabled));
NEMR4T g357(.s(next_interrupt_enabled1), .d(next_interrupt_enabled10), .b(vdd), .g(inst[0]));
NEMR4T g358(.s(next_interrupt_enabled10), .d(AA_345), .b(vdd), .g(inst[16]));
NEMR4T g359(.s(AA_345), .d(AA_344), .b(vdd), .g(inst[13]));
NEMR4T g360(.s(AA_344), .d(AA_360), .b(vdd), .g(irq));
NEMR4T g361(.s(AA_344), .d(AA_397), .b(gnd), .g(irq));
NEMR4T g362(.s(AA_345), .d(AA_344), .b(gnd), .g(inst[13]));
NEMR4T g363(.s(next_interrupt_enabled10), .d(next_interrupt_enabled101), .b(gnd), .g(inst[16]));
NEMR4T g364(.s(next_interrupt_enabled101), .d(next_interrupt_enabled1010), .b(vdd), .g(inst[13]));
NEMR4T g365(.s(next_interrupt_enabled1010), .d(next_interrupt_enabled10100), .b(vdd), .g(irq));
NEMR4T g366(.s(next_interrupt_enabled10100), .d(AA_388), .b(vdd), .g(inst[17]));
NEMR4T g367(.s(next_interrupt_enabled10100), .d(AA_382), .b(gnd), .g(inst[17]));
NEMR4T g368(.s(next_interrupt_enabled1010), .d(AA_397), .b(gnd), .g(irq));
NEMR4T g369(.s(next_interrupt_enabled101), .d(AA_344), .b(gnd), .g(inst[13]));
NEMR4T g370(.s(next_interrupt_enabled1), .d(next_interrupt_enabled11), .b(gnd), .g(inst[0]));
NEMR4T g371(.s(next_interrupt_enabled11), .d(AA_345), .b(vdd), .g(inst[16]));
NEMR4T g372(.s(next_interrupt_enabled11), .d(AA_345), .b(gnd), .g(inst[16]));
NEMR4T g373(.s(werf), .d(werf0), .b(vdd), .g(inst[14]));
NEMR4T g374(.s(werf0), .d(werf00), .b(vdd), .g(inst[16]));
NEMR4T g375(.s(werf00), .d(werf000), .b(vdd), .g(inst[13]));
NEMR4T g376(.s(werf000), .d(werf0000), .b(vdd), .g(irq));
NEMR4T g377(.s(werf0000), .d(AA_382), .b(vdd), .g(inst[17]));
NEMR4T g378(.s(werf0000), .d(AA_382), .b(gnd), .g(inst[17]));
NEMR4T g379(.s(werf000), .d(AA_397), .b(gnd), .g(irq));
NEMR4T g380(.s(werf00), .d(AA_386), .b(gnd), .g(inst[13]));
NEMR4T g381(.s(werf0), .d(AA_387), .b(gnd), .g(inst[16]));
NEMR4T g382(.s(werf), .d(werf1), .b(gnd), .g(inst[14]));
NEMR4T g383(.s(werf1), .d(werf10), .b(vdd), .g(inst[16]));
NEMR4T g384(.s(werf10), .d(AA_375), .b(vdd), .g(inst[13]));
NEMR4T g385(.s(AA_375), .d(AA_374), .b(vdd), .g(irq));
NEMR4T g386(.s(AA_374), .d(AA_388), .b(vdd), .g(inst[17]));
NEMR4T g387(.s(AA_374), .d(AA_396), .b(gnd), .g(inst[17]));
NEMR4T g388(.s(AA_375), .d(AA_397), .b(gnd), .g(irq));
NEMR4T g389(.s(werf10), .d(AA_375), .b(gnd), .g(inst[13]));
NEMR4T g390(.s(werf1), .d(AA_387), .b(gnd), .g(inst[16]));
NEMR4T g391(.s(wesp), .d(AA_403), .b(vdd), .g(inst[14]));
NEMR4T g392(.s(wesp), .d(wesp1), .b(gnd), .g(inst[14]));
NEMR4T g393(.s(wesp1), .d(AA_404), .b(vdd), .g(inst[16]));
NEMR4T g394(.s(wesp1), .d(AA_400), .b(gnd), .g(inst[16]));

endmodule